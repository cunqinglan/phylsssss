module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 ;
  wire n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n341 , n342 , n343 , n345 , n346 , n347 , n348 , n349 , n350 , n352 , n353 , n354 , n355 , n356 , n358 , n359 , n360 , n361 , n362 , n364 , n365 , n367 , n368 , n369 , n370 , n371 , n373 , n374 , n375 , n376 , n377 , n379 , n380 , n382 , n383 , n384 , n385 , n386 , n388 , n389 , n390 , n391 , n392 , n394 , n395 , n397 , n398 , n399 , n400 , n401 , n403 , n404 , n405 , n406 , n407 , n409 , n410 , n412 , n413 , n414 , n415 , n416 , n418 , n419 , n420 , n421 , n422 , n424 , n425 , n427 , n428 , n429 , n430 , n431 , n433 , n434 , n435 , n436 , n437 , n439 , n440 , n442 , n443 , n444 , n445 , n446 , n448 , n449 , n450 , n451 , n452 , n454 , n455 , n457 , n458 , n459 , n460 , n461 , n463 , n464 , n465 , n466 , n467 , n469 , n470 , n472 , n473 , n474 , n475 , n476 , n478 , n479 , n480 , n481 , n482 , n484 , n485 , n487 , n488 , n489 , n490 , n491 , n493 , n494 , n495 , n496 , n497 , n499 , n500 , n502 , n503 , n504 , n505 , n506 , n508 , n509 , n510 , n511 , n512 , n514 , n515 , n517 , n518 , n519 , n520 , n521 , n523 , n524 , n525 , n526 , n527 , n529 , n530 , n532 , n533 , n534 , n535 , n536 , n538 , n539 , n540 , n541 , n542 , n544 , n545 , n547 , n548 , n549 , n550 , n551 , n553 , n554 , n555 , n556 , n557 , n559 , n560 , n562 , n563 , n564 , n565 , n566 , n568 , n569 , n570 , n571 , n572 , n574 , n575 , n577 , n578 , n579 , n580 , n581 , n583 , n584 , n585 , n586 , n587 , n589 , n590 , n592 , n593 , n594 , n595 , n596 , n598 , n599 , n600 , n601 , n602 , n604 , n605 , n607 , n608 , n609 , n610 , n611 , n613 , n614 , n615 , n616 , n617 , n619 , n620 , n622 , n623 , n624 , n625 , n626 , n628 , n629 , n630 , n631 , n632 , n634 , n635 , n637 , n638 , n639 , n640 , n641 , n643 , n644 , n645 , n646 , n647 , n649 , n650 , n652 , n653 , n654 , n655 , n656 , n658 , n659 , n660 , n661 , n662 , n664 , n665 , n667 , n668 , n669 , n670 , n671 , n673 , n674 , n675 , n676 , n677 , n679 , n680 , n682 , n683 , n684 , n685 , n686 , n688 , n689 , n690 , n691 , n692 , n694 , n695 , n697 , n698 , n699 , n700 , n701 , n703 , n704 , n705 , n706 , n707 , n709 , n710 , n712 , n713 , n714 , n715 , n716 , n718 , n719 , n720 , n721 , n722 , n724 , n725 , n727 , n728 , n729 , n730 , n731 , n733 , n734 , n735 , n736 , n737 , n739 , n740 , n742 , n743 , n744 , n745 , n746 , n748 , n749 , n750 , n751 , n752 , n754 , n755 , n757 , n758 , n759 , n760 , n761 , n763 , n764 , n765 , n766 , n767 , n769 , n770 , n772 , n773 , n774 , n775 , n776 , n778 , n779 , n780 , n781 , n782 , n784 , n785 , n787 , n788 , n789 , n790 , n791 , n793 , n794 , n795 , n796 , n797 , n799 , n800 , n802 , n803 , n804 , n805 , n806 , n808 , n809 , n810 , n811 , n812 , n814 , n815 , n817 , n818 , n819 , n820 , n821 , n823 , n824 , n825 , n826 , n827 , n829 , n830 , n832 , n833 , n834 , n835 , n836 , n838 , n839 , n840 , n841 , n842 , n844 , n845 , n847 , n848 , n849 , n850 , n851 , n853 , n854 , n855 , n856 , n857 , n859 , n860 , n862 , n863 , n864 , n865 , n866 , n868 , n869 , n870 , n871 , n872 , n874 , n875 , n877 , n878 , n879 , n880 , n881 , n883 , n884 , n885 , n886 , n887 , n889 , n890 , n892 , n893 , n894 , n895 , n896 , n898 , n899 , n900 , n901 , n902 , n904 , n905 , n907 , n908 , n909 , n910 , n911 , n913 , n914 , n915 , n916 , n917 , n919 , n920 , n922 , n923 , n924 , n925 , n926 , n928 , n929 , n930 , n931 , n932 , n934 , n935 , n937 , n938 , n939 , n940 , n941 , n943 , n944 , n945 , n946 , n947 , n949 , n950 , n952 , n953 , n954 , n955 , n956 , n958 , n959 , n960 , n961 , n962 , n964 , n965 , n967 , n968 , n969 , n970 , n972 , n973 , n974 , n975 , n976 ;
  XOR2xp5_ASAP7_75t_R       g000( .A (x0), .B (x128), .Y (y0) );
  NAND2xp33_ASAP7_75t_R     g001( .A (x0), .B (x128), .Y (n341) );
  XNOR2xp5_ASAP7_75t_R      g002( .A (x1), .B (x129), .Y (n343) );
  XOR2xp5_ASAP7_75t_R       g003( .A (n341), .B (n343), .Y (y1) );
  NAND2xp33_ASAP7_75t_R     g004( .A (x1), .B (x129), .Y (n342) );
  OAI211xp5_ASAP7_75t_R     g005( .A1 (x1), .A2 (x129), .B (x128), .C (x0), .Y (n345) );
  NAND2xp33_ASAP7_75t_R     g006( .A (n342), .B (n345), .Y (n346) );
  NOR2xp33_ASAP7_75t_R      g007( .A (x2), .B (x130), .Y (n347) );
  NAND2xp33_ASAP7_75t_R     g008( .A (x2), .B (x130), .Y (n348) );
  INVx1_ASAP7_75t_R         g009( .A (n348), .Y (n349) );
  NOR2xp33_ASAP7_75t_R      g010( .A (n347), .B (n349), .Y (n350) );
  XOR2xp5_ASAP7_75t_R       g011( .A (n346), .B (n350), .Y (y2) );
  A2O1A1Ixp33_ASAP7_75t_R   g012( .A1 (n342), .B (n347), .A2 (n345), .C (n348), .Y (n352) );
  NOR2xp33_ASAP7_75t_R      g013( .A (x3), .B (x131), .Y (n353) );
  AND2x2_ASAP7_75t_R        g014( .A (x3), .B (x131), .Y (n355) );
  NOR2xp33_ASAP7_75t_R      g015( .A (n353), .B (n355), .Y (n356) );
  XOR2xp5_ASAP7_75t_R       g016( .A (n352), .B (n356), .Y (y3) );
  OR2x2_ASAP7_75t_R         g017( .A (x4), .B (x132), .Y (n359) );
  NAND2xp33_ASAP7_75t_R     g018( .A (x4), .B (x132), .Y (n360) );
  NAND2xp33_ASAP7_75t_R     g019( .A (n359), .B (n360), .Y (n362) );
  INVx1_ASAP7_75t_R         g020( .A (n353), .Y (n354) );
  AOI21xp33_ASAP7_75t_R     g021( .A1 (n352), .B (n355), .A2 (n354), .Y (n358) );
  XOR2xp5_ASAP7_75t_R       g022( .A (n362), .B (n358), .Y (y4) );
  XNOR2xp5_ASAP7_75t_R      g023( .A (x5), .B (x133), .Y (n365) );
  INVx1_ASAP7_75t_R         g024( .A (n360), .Y (n361) );
  A2O1A1O1Ixp25_ASAP7_75t_R g025( .A1 (n352), .B (n355), .D (n361), .A2 (n354), .C (n359), .Y (n364) );
  XOR2xp5_ASAP7_75t_R       g026( .A (n365), .B (n364), .Y (y5) );
  INVx1_ASAP7_75t_R         g027( .A (x5), .Y (n258) );
  INVx1_ASAP7_75t_R         g028( .A (x133), .Y (n299) );
  MAJIxp5_ASAP7_75t_R       g029( .A (n258), .B (n299), .C (n364), .Y (n367) );
  NOR2xp33_ASAP7_75t_R      g030( .A (x6), .B (x134), .Y (n368) );
  AND2x2_ASAP7_75t_R        g031( .A (x6), .B (x134), .Y (n370) );
  NOR2xp33_ASAP7_75t_R      g032( .A (n368), .B (n370), .Y (n371) );
  XOR2xp5_ASAP7_75t_R       g033( .A (n367), .B (n371), .Y (y6) );
  OR2x2_ASAP7_75t_R         g034( .A (x7), .B (x135), .Y (n374) );
  NAND2xp33_ASAP7_75t_R     g035( .A (x7), .B (x135), .Y (n375) );
  NAND2xp33_ASAP7_75t_R     g036( .A (n374), .B (n375), .Y (n377) );
  INVx1_ASAP7_75t_R         g037( .A (n368), .Y (n369) );
  AOI21xp33_ASAP7_75t_R     g038( .A1 (n367), .B (n370), .A2 (n369), .Y (n373) );
  XOR2xp5_ASAP7_75t_R       g039( .A (n377), .B (n373), .Y (y7) );
  XNOR2xp5_ASAP7_75t_R      g040( .A (x8), .B (x136), .Y (n380) );
  INVx1_ASAP7_75t_R         g041( .A (n375), .Y (n376) );
  A2O1A1O1Ixp25_ASAP7_75t_R g042( .A1 (n367), .B (n370), .D (n376), .A2 (n369), .C (n374), .Y (n379) );
  XOR2xp5_ASAP7_75t_R       g043( .A (n380), .B (n379), .Y (y8) );
  INVx1_ASAP7_75t_R         g044( .A (x8), .Y (n259) );
  INVx1_ASAP7_75t_R         g045( .A (x136), .Y (n300) );
  MAJIxp5_ASAP7_75t_R       g046( .A (n259), .B (n300), .C (n379), .Y (n382) );
  NOR2xp33_ASAP7_75t_R      g047( .A (x9), .B (x137), .Y (n383) );
  AND2x2_ASAP7_75t_R        g048( .A (x9), .B (x137), .Y (n385) );
  NOR2xp33_ASAP7_75t_R      g049( .A (n383), .B (n385), .Y (n386) );
  XOR2xp5_ASAP7_75t_R       g050( .A (n382), .B (n386), .Y (y9) );
  OR2x2_ASAP7_75t_R         g051( .A (x10), .B (x138), .Y (n389) );
  NAND2xp33_ASAP7_75t_R     g052( .A (x10), .B (x138), .Y (n390) );
  NAND2xp33_ASAP7_75t_R     g053( .A (n389), .B (n390), .Y (n392) );
  INVx1_ASAP7_75t_R         g054( .A (n383), .Y (n384) );
  AOI21xp33_ASAP7_75t_R     g055( .A1 (n382), .B (n385), .A2 (n384), .Y (n388) );
  XOR2xp5_ASAP7_75t_R       g056( .A (n392), .B (n388), .Y (y10) );
  XNOR2xp5_ASAP7_75t_R      g057( .A (x11), .B (x139), .Y (n395) );
  INVx1_ASAP7_75t_R         g058( .A (n390), .Y (n391) );
  A2O1A1O1Ixp25_ASAP7_75t_R g059( .A1 (n382), .B (n385), .D (n391), .A2 (n384), .C (n389), .Y (n394) );
  XOR2xp5_ASAP7_75t_R       g060( .A (n395), .B (n394), .Y (y11) );
  INVx1_ASAP7_75t_R         g061( .A (x11), .Y (n260) );
  INVx1_ASAP7_75t_R         g062( .A (x139), .Y (n301) );
  MAJIxp5_ASAP7_75t_R       g063( .A (n260), .B (n301), .C (n394), .Y (n397) );
  NOR2xp33_ASAP7_75t_R      g064( .A (x12), .B (x140), .Y (n398) );
  AND2x2_ASAP7_75t_R        g065( .A (x12), .B (x140), .Y (n400) );
  NOR2xp33_ASAP7_75t_R      g066( .A (n398), .B (n400), .Y (n401) );
  XOR2xp5_ASAP7_75t_R       g067( .A (n397), .B (n401), .Y (y12) );
  OR2x2_ASAP7_75t_R         g068( .A (x13), .B (x141), .Y (n404) );
  NAND2xp33_ASAP7_75t_R     g069( .A (x13), .B (x141), .Y (n405) );
  NAND2xp33_ASAP7_75t_R     g070( .A (n404), .B (n405), .Y (n407) );
  INVx1_ASAP7_75t_R         g071( .A (n398), .Y (n399) );
  AOI21xp33_ASAP7_75t_R     g072( .A1 (n397), .B (n400), .A2 (n399), .Y (n403) );
  XOR2xp5_ASAP7_75t_R       g073( .A (n407), .B (n403), .Y (y13) );
  XNOR2xp5_ASAP7_75t_R      g074( .A (x14), .B (x142), .Y (n410) );
  INVx1_ASAP7_75t_R         g075( .A (n405), .Y (n406) );
  A2O1A1O1Ixp25_ASAP7_75t_R g076( .A1 (n397), .B (n400), .D (n406), .A2 (n399), .C (n404), .Y (n409) );
  XOR2xp5_ASAP7_75t_R       g077( .A (n410), .B (n409), .Y (y14) );
  INVx1_ASAP7_75t_R         g078( .A (x14), .Y (n261) );
  INVx1_ASAP7_75t_R         g079( .A (x142), .Y (n302) );
  MAJIxp5_ASAP7_75t_R       g080( .A (n261), .B (n302), .C (n409), .Y (n412) );
  NOR2xp33_ASAP7_75t_R      g081( .A (x15), .B (x143), .Y (n413) );
  AND2x2_ASAP7_75t_R        g082( .A (x15), .B (x143), .Y (n415) );
  NOR2xp33_ASAP7_75t_R      g083( .A (n413), .B (n415), .Y (n416) );
  XOR2xp5_ASAP7_75t_R       g084( .A (n412), .B (n416), .Y (y15) );
  OR2x2_ASAP7_75t_R         g085( .A (x16), .B (x144), .Y (n419) );
  NAND2xp33_ASAP7_75t_R     g086( .A (x16), .B (x144), .Y (n420) );
  NAND2xp33_ASAP7_75t_R     g087( .A (n419), .B (n420), .Y (n422) );
  INVx1_ASAP7_75t_R         g088( .A (n413), .Y (n414) );
  AOI21xp33_ASAP7_75t_R     g089( .A1 (n412), .B (n415), .A2 (n414), .Y (n418) );
  XOR2xp5_ASAP7_75t_R       g090( .A (n422), .B (n418), .Y (y16) );
  XNOR2xp5_ASAP7_75t_R      g091( .A (x17), .B (x145), .Y (n425) );
  INVx1_ASAP7_75t_R         g092( .A (n420), .Y (n421) );
  A2O1A1O1Ixp25_ASAP7_75t_R g093( .A1 (n412), .B (n415), .D (n421), .A2 (n414), .C (n419), .Y (n424) );
  XOR2xp5_ASAP7_75t_R       g094( .A (n425), .B (n424), .Y (y17) );
  INVx1_ASAP7_75t_R         g095( .A (x17), .Y (n262) );
  INVx1_ASAP7_75t_R         g096( .A (x145), .Y (n303) );
  MAJIxp5_ASAP7_75t_R       g097( .A (n262), .B (n303), .C (n424), .Y (n427) );
  NOR2xp33_ASAP7_75t_R      g098( .A (x18), .B (x146), .Y (n428) );
  AND2x2_ASAP7_75t_R        g099( .A (x18), .B (x146), .Y (n430) );
  NOR2xp33_ASAP7_75t_R      g100( .A (n428), .B (n430), .Y (n431) );
  XOR2xp5_ASAP7_75t_R       g101( .A (n427), .B (n431), .Y (y18) );
  OR2x2_ASAP7_75t_R         g102( .A (x19), .B (x147), .Y (n434) );
  NAND2xp33_ASAP7_75t_R     g103( .A (x19), .B (x147), .Y (n435) );
  NAND2xp33_ASAP7_75t_R     g104( .A (n434), .B (n435), .Y (n437) );
  INVx1_ASAP7_75t_R         g105( .A (n428), .Y (n429) );
  AOI21xp33_ASAP7_75t_R     g106( .A1 (n427), .B (n430), .A2 (n429), .Y (n433) );
  XOR2xp5_ASAP7_75t_R       g107( .A (n437), .B (n433), .Y (y19) );
  XNOR2xp5_ASAP7_75t_R      g108( .A (x20), .B (x148), .Y (n440) );
  INVx1_ASAP7_75t_R         g109( .A (n435), .Y (n436) );
  A2O1A1O1Ixp25_ASAP7_75t_R g110( .A1 (n427), .B (n430), .D (n436), .A2 (n429), .C (n434), .Y (n439) );
  XOR2xp5_ASAP7_75t_R       g111( .A (n440), .B (n439), .Y (y20) );
  INVx1_ASAP7_75t_R         g112( .A (x20), .Y (n263) );
  INVx1_ASAP7_75t_R         g113( .A (x148), .Y (n304) );
  MAJIxp5_ASAP7_75t_R       g114( .A (n263), .B (n304), .C (n439), .Y (n442) );
  NOR2xp33_ASAP7_75t_R      g115( .A (x21), .B (x149), .Y (n443) );
  AND2x2_ASAP7_75t_R        g116( .A (x21), .B (x149), .Y (n445) );
  NOR2xp33_ASAP7_75t_R      g117( .A (n443), .B (n445), .Y (n446) );
  XOR2xp5_ASAP7_75t_R       g118( .A (n442), .B (n446), .Y (y21) );
  OR2x2_ASAP7_75t_R         g119( .A (x22), .B (x150), .Y (n449) );
  NAND2xp33_ASAP7_75t_R     g120( .A (x22), .B (x150), .Y (n450) );
  NAND2xp33_ASAP7_75t_R     g121( .A (n449), .B (n450), .Y (n452) );
  INVx1_ASAP7_75t_R         g122( .A (n443), .Y (n444) );
  AOI21xp33_ASAP7_75t_R     g123( .A1 (n442), .B (n445), .A2 (n444), .Y (n448) );
  XOR2xp5_ASAP7_75t_R       g124( .A (n452), .B (n448), .Y (y22) );
  XNOR2xp5_ASAP7_75t_R      g125( .A (x23), .B (x151), .Y (n455) );
  INVx1_ASAP7_75t_R         g126( .A (n450), .Y (n451) );
  A2O1A1O1Ixp25_ASAP7_75t_R g127( .A1 (n442), .B (n445), .D (n451), .A2 (n444), .C (n449), .Y (n454) );
  XOR2xp5_ASAP7_75t_R       g128( .A (n455), .B (n454), .Y (y23) );
  INVx1_ASAP7_75t_R         g129( .A (x23), .Y (n264) );
  INVx1_ASAP7_75t_R         g130( .A (x151), .Y (n305) );
  MAJIxp5_ASAP7_75t_R       g131( .A (n264), .B (n305), .C (n454), .Y (n457) );
  NOR2xp33_ASAP7_75t_R      g132( .A (x24), .B (x152), .Y (n458) );
  AND2x2_ASAP7_75t_R        g133( .A (x24), .B (x152), .Y (n460) );
  NOR2xp33_ASAP7_75t_R      g134( .A (n458), .B (n460), .Y (n461) );
  XOR2xp5_ASAP7_75t_R       g135( .A (n457), .B (n461), .Y (y24) );
  OR2x2_ASAP7_75t_R         g136( .A (x25), .B (x153), .Y (n464) );
  NAND2xp33_ASAP7_75t_R     g137( .A (x25), .B (x153), .Y (n465) );
  NAND2xp33_ASAP7_75t_R     g138( .A (n464), .B (n465), .Y (n467) );
  INVx1_ASAP7_75t_R         g139( .A (n458), .Y (n459) );
  AOI21xp33_ASAP7_75t_R     g140( .A1 (n457), .B (n460), .A2 (n459), .Y (n463) );
  XOR2xp5_ASAP7_75t_R       g141( .A (n467), .B (n463), .Y (y25) );
  XNOR2xp5_ASAP7_75t_R      g142( .A (x26), .B (x154), .Y (n470) );
  INVx1_ASAP7_75t_R         g143( .A (n465), .Y (n466) );
  A2O1A1O1Ixp25_ASAP7_75t_R g144( .A1 (n457), .B (n460), .D (n466), .A2 (n459), .C (n464), .Y (n469) );
  XOR2xp5_ASAP7_75t_R       g145( .A (n470), .B (n469), .Y (y26) );
  INVx1_ASAP7_75t_R         g146( .A (x26), .Y (n265) );
  INVx1_ASAP7_75t_R         g147( .A (x154), .Y (n306) );
  MAJIxp5_ASAP7_75t_R       g148( .A (n265), .B (n306), .C (n469), .Y (n472) );
  NOR2xp33_ASAP7_75t_R      g149( .A (x27), .B (x155), .Y (n473) );
  AND2x2_ASAP7_75t_R        g150( .A (x27), .B (x155), .Y (n475) );
  NOR2xp33_ASAP7_75t_R      g151( .A (n473), .B (n475), .Y (n476) );
  XOR2xp5_ASAP7_75t_R       g152( .A (n472), .B (n476), .Y (y27) );
  OR2x2_ASAP7_75t_R         g153( .A (x28), .B (x156), .Y (n479) );
  NAND2xp33_ASAP7_75t_R     g154( .A (x28), .B (x156), .Y (n480) );
  NAND2xp33_ASAP7_75t_R     g155( .A (n479), .B (n480), .Y (n482) );
  INVx1_ASAP7_75t_R         g156( .A (n473), .Y (n474) );
  AOI21xp33_ASAP7_75t_R     g157( .A1 (n472), .B (n475), .A2 (n474), .Y (n478) );
  XOR2xp5_ASAP7_75t_R       g158( .A (n482), .B (n478), .Y (y28) );
  XNOR2xp5_ASAP7_75t_R      g159( .A (x29), .B (x157), .Y (n485) );
  INVx1_ASAP7_75t_R         g160( .A (n480), .Y (n481) );
  A2O1A1O1Ixp25_ASAP7_75t_R g161( .A1 (n472), .B (n475), .D (n481), .A2 (n474), .C (n479), .Y (n484) );
  XOR2xp5_ASAP7_75t_R       g162( .A (n485), .B (n484), .Y (y29) );
  INVx1_ASAP7_75t_R         g163( .A (x29), .Y (n266) );
  INVx1_ASAP7_75t_R         g164( .A (x157), .Y (n307) );
  MAJIxp5_ASAP7_75t_R       g165( .A (n266), .B (n307), .C (n484), .Y (n487) );
  NOR2xp33_ASAP7_75t_R      g166( .A (x30), .B (x158), .Y (n488) );
  AND2x2_ASAP7_75t_R        g167( .A (x30), .B (x158), .Y (n490) );
  NOR2xp33_ASAP7_75t_R      g168( .A (n488), .B (n490), .Y (n491) );
  XOR2xp5_ASAP7_75t_R       g169( .A (n487), .B (n491), .Y (y30) );
  OR2x2_ASAP7_75t_R         g170( .A (x31), .B (x159), .Y (n494) );
  NAND2xp33_ASAP7_75t_R     g171( .A (x31), .B (x159), .Y (n495) );
  NAND2xp33_ASAP7_75t_R     g172( .A (n494), .B (n495), .Y (n497) );
  INVx1_ASAP7_75t_R         g173( .A (n488), .Y (n489) );
  AOI21xp33_ASAP7_75t_R     g174( .A1 (n487), .B (n490), .A2 (n489), .Y (n493) );
  XOR2xp5_ASAP7_75t_R       g175( .A (n497), .B (n493), .Y (y31) );
  XNOR2xp5_ASAP7_75t_R      g176( .A (x32), .B (x160), .Y (n500) );
  INVx1_ASAP7_75t_R         g177( .A (n495), .Y (n496) );
  A2O1A1O1Ixp25_ASAP7_75t_R g178( .A1 (n487), .B (n490), .D (n496), .A2 (n489), .C (n494), .Y (n499) );
  XOR2xp5_ASAP7_75t_R       g179( .A (n500), .B (n499), .Y (y32) );
  INVx1_ASAP7_75t_R         g180( .A (x32), .Y (n267) );
  INVx1_ASAP7_75t_R         g181( .A (x160), .Y (n308) );
  MAJIxp5_ASAP7_75t_R       g182( .A (n267), .B (n308), .C (n499), .Y (n502) );
  NOR2xp33_ASAP7_75t_R      g183( .A (x33), .B (x161), .Y (n503) );
  AND2x2_ASAP7_75t_R        g184( .A (x33), .B (x161), .Y (n505) );
  NOR2xp33_ASAP7_75t_R      g185( .A (n503), .B (n505), .Y (n506) );
  XOR2xp5_ASAP7_75t_R       g186( .A (n502), .B (n506), .Y (y33) );
  OR2x2_ASAP7_75t_R         g187( .A (x34), .B (x162), .Y (n509) );
  NAND2xp33_ASAP7_75t_R     g188( .A (x34), .B (x162), .Y (n510) );
  NAND2xp33_ASAP7_75t_R     g189( .A (n509), .B (n510), .Y (n512) );
  INVx1_ASAP7_75t_R         g190( .A (n503), .Y (n504) );
  AOI21xp33_ASAP7_75t_R     g191( .A1 (n502), .B (n505), .A2 (n504), .Y (n508) );
  XOR2xp5_ASAP7_75t_R       g192( .A (n512), .B (n508), .Y (y34) );
  XNOR2xp5_ASAP7_75t_R      g193( .A (x35), .B (x163), .Y (n515) );
  INVx1_ASAP7_75t_R         g194( .A (n510), .Y (n511) );
  A2O1A1O1Ixp25_ASAP7_75t_R g195( .A1 (n502), .B (n505), .D (n511), .A2 (n504), .C (n509), .Y (n514) );
  XOR2xp5_ASAP7_75t_R       g196( .A (n515), .B (n514), .Y (y35) );
  INVx1_ASAP7_75t_R         g197( .A (x35), .Y (n268) );
  INVx1_ASAP7_75t_R         g198( .A (x163), .Y (n309) );
  MAJIxp5_ASAP7_75t_R       g199( .A (n268), .B (n309), .C (n514), .Y (n517) );
  NOR2xp33_ASAP7_75t_R      g200( .A (x36), .B (x164), .Y (n518) );
  AND2x2_ASAP7_75t_R        g201( .A (x36), .B (x164), .Y (n520) );
  NOR2xp33_ASAP7_75t_R      g202( .A (n518), .B (n520), .Y (n521) );
  XOR2xp5_ASAP7_75t_R       g203( .A (n517), .B (n521), .Y (y36) );
  OR2x2_ASAP7_75t_R         g204( .A (x37), .B (x165), .Y (n524) );
  NAND2xp33_ASAP7_75t_R     g205( .A (x37), .B (x165), .Y (n525) );
  NAND2xp33_ASAP7_75t_R     g206( .A (n524), .B (n525), .Y (n527) );
  INVx1_ASAP7_75t_R         g207( .A (n518), .Y (n519) );
  AOI21xp33_ASAP7_75t_R     g208( .A1 (n517), .B (n520), .A2 (n519), .Y (n523) );
  XOR2xp5_ASAP7_75t_R       g209( .A (n527), .B (n523), .Y (y37) );
  XNOR2xp5_ASAP7_75t_R      g210( .A (x38), .B (x166), .Y (n530) );
  INVx1_ASAP7_75t_R         g211( .A (n525), .Y (n526) );
  A2O1A1O1Ixp25_ASAP7_75t_R g212( .A1 (n517), .B (n520), .D (n526), .A2 (n519), .C (n524), .Y (n529) );
  XOR2xp5_ASAP7_75t_R       g213( .A (n530), .B (n529), .Y (y38) );
  INVx1_ASAP7_75t_R         g214( .A (x38), .Y (n269) );
  INVx1_ASAP7_75t_R         g215( .A (x166), .Y (n310) );
  MAJIxp5_ASAP7_75t_R       g216( .A (n269), .B (n310), .C (n529), .Y (n532) );
  NOR2xp33_ASAP7_75t_R      g217( .A (x39), .B (x167), .Y (n533) );
  AND2x2_ASAP7_75t_R        g218( .A (x39), .B (x167), .Y (n535) );
  NOR2xp33_ASAP7_75t_R      g219( .A (n533), .B (n535), .Y (n536) );
  XOR2xp5_ASAP7_75t_R       g220( .A (n532), .B (n536), .Y (y39) );
  OR2x2_ASAP7_75t_R         g221( .A (x40), .B (x168), .Y (n539) );
  NAND2xp33_ASAP7_75t_R     g222( .A (x40), .B (x168), .Y (n540) );
  NAND2xp33_ASAP7_75t_R     g223( .A (n539), .B (n540), .Y (n542) );
  INVx1_ASAP7_75t_R         g224( .A (n533), .Y (n534) );
  AOI21xp33_ASAP7_75t_R     g225( .A1 (n532), .B (n535), .A2 (n534), .Y (n538) );
  XOR2xp5_ASAP7_75t_R       g226( .A (n542), .B (n538), .Y (y40) );
  XNOR2xp5_ASAP7_75t_R      g227( .A (x41), .B (x169), .Y (n545) );
  INVx1_ASAP7_75t_R         g228( .A (n540), .Y (n541) );
  A2O1A1O1Ixp25_ASAP7_75t_R g229( .A1 (n532), .B (n535), .D (n541), .A2 (n534), .C (n539), .Y (n544) );
  XOR2xp5_ASAP7_75t_R       g230( .A (n545), .B (n544), .Y (y41) );
  INVx1_ASAP7_75t_R         g231( .A (x41), .Y (n270) );
  INVx1_ASAP7_75t_R         g232( .A (x169), .Y (n311) );
  MAJIxp5_ASAP7_75t_R       g233( .A (n270), .B (n311), .C (n544), .Y (n547) );
  NOR2xp33_ASAP7_75t_R      g234( .A (x42), .B (x170), .Y (n548) );
  AND2x2_ASAP7_75t_R        g235( .A (x42), .B (x170), .Y (n550) );
  NOR2xp33_ASAP7_75t_R      g236( .A (n548), .B (n550), .Y (n551) );
  XOR2xp5_ASAP7_75t_R       g237( .A (n547), .B (n551), .Y (y42) );
  OR2x2_ASAP7_75t_R         g238( .A (x43), .B (x171), .Y (n554) );
  NAND2xp33_ASAP7_75t_R     g239( .A (x43), .B (x171), .Y (n555) );
  NAND2xp33_ASAP7_75t_R     g240( .A (n554), .B (n555), .Y (n557) );
  INVx1_ASAP7_75t_R         g241( .A (n548), .Y (n549) );
  AOI21xp33_ASAP7_75t_R     g242( .A1 (n547), .B (n550), .A2 (n549), .Y (n553) );
  XOR2xp5_ASAP7_75t_R       g243( .A (n557), .B (n553), .Y (y43) );
  XNOR2xp5_ASAP7_75t_R      g244( .A (x44), .B (x172), .Y (n560) );
  INVx1_ASAP7_75t_R         g245( .A (n555), .Y (n556) );
  A2O1A1O1Ixp25_ASAP7_75t_R g246( .A1 (n547), .B (n550), .D (n556), .A2 (n549), .C (n554), .Y (n559) );
  XOR2xp5_ASAP7_75t_R       g247( .A (n560), .B (n559), .Y (y44) );
  INVx1_ASAP7_75t_R         g248( .A (x44), .Y (n271) );
  INVx1_ASAP7_75t_R         g249( .A (x172), .Y (n312) );
  MAJIxp5_ASAP7_75t_R       g250( .A (n271), .B (n312), .C (n559), .Y (n562) );
  NOR2xp33_ASAP7_75t_R      g251( .A (x45), .B (x173), .Y (n563) );
  AND2x2_ASAP7_75t_R        g252( .A (x45), .B (x173), .Y (n565) );
  NOR2xp33_ASAP7_75t_R      g253( .A (n563), .B (n565), .Y (n566) );
  XOR2xp5_ASAP7_75t_R       g254( .A (n562), .B (n566), .Y (y45) );
  OR2x2_ASAP7_75t_R         g255( .A (x46), .B (x174), .Y (n569) );
  NAND2xp33_ASAP7_75t_R     g256( .A (x46), .B (x174), .Y (n570) );
  NAND2xp33_ASAP7_75t_R     g257( .A (n569), .B (n570), .Y (n572) );
  INVx1_ASAP7_75t_R         g258( .A (n563), .Y (n564) );
  AOI21xp33_ASAP7_75t_R     g259( .A1 (n562), .B (n565), .A2 (n564), .Y (n568) );
  XOR2xp5_ASAP7_75t_R       g260( .A (n572), .B (n568), .Y (y46) );
  XNOR2xp5_ASAP7_75t_R      g261( .A (x47), .B (x175), .Y (n575) );
  INVx1_ASAP7_75t_R         g262( .A (n570), .Y (n571) );
  A2O1A1O1Ixp25_ASAP7_75t_R g263( .A1 (n562), .B (n565), .D (n571), .A2 (n564), .C (n569), .Y (n574) );
  XOR2xp5_ASAP7_75t_R       g264( .A (n575), .B (n574), .Y (y47) );
  INVx1_ASAP7_75t_R         g265( .A (x47), .Y (n272) );
  INVx1_ASAP7_75t_R         g266( .A (x175), .Y (n313) );
  MAJIxp5_ASAP7_75t_R       g267( .A (n272), .B (n313), .C (n574), .Y (n577) );
  NOR2xp33_ASAP7_75t_R      g268( .A (x48), .B (x176), .Y (n578) );
  AND2x2_ASAP7_75t_R        g269( .A (x48), .B (x176), .Y (n580) );
  NOR2xp33_ASAP7_75t_R      g270( .A (n578), .B (n580), .Y (n581) );
  XOR2xp5_ASAP7_75t_R       g271( .A (n577), .B (n581), .Y (y48) );
  OR2x2_ASAP7_75t_R         g272( .A (x49), .B (x177), .Y (n584) );
  NAND2xp33_ASAP7_75t_R     g273( .A (x49), .B (x177), .Y (n585) );
  NAND2xp33_ASAP7_75t_R     g274( .A (n584), .B (n585), .Y (n587) );
  INVx1_ASAP7_75t_R         g275( .A (n578), .Y (n579) );
  AOI21xp33_ASAP7_75t_R     g276( .A1 (n577), .B (n580), .A2 (n579), .Y (n583) );
  XOR2xp5_ASAP7_75t_R       g277( .A (n587), .B (n583), .Y (y49) );
  XNOR2xp5_ASAP7_75t_R      g278( .A (x50), .B (x178), .Y (n590) );
  INVx1_ASAP7_75t_R         g279( .A (n585), .Y (n586) );
  A2O1A1O1Ixp25_ASAP7_75t_R g280( .A1 (n577), .B (n580), .D (n586), .A2 (n579), .C (n584), .Y (n589) );
  XOR2xp5_ASAP7_75t_R       g281( .A (n590), .B (n589), .Y (y50) );
  INVx1_ASAP7_75t_R         g282( .A (x50), .Y (n273) );
  INVx1_ASAP7_75t_R         g283( .A (x178), .Y (n314) );
  MAJIxp5_ASAP7_75t_R       g284( .A (n273), .B (n314), .C (n589), .Y (n592) );
  NOR2xp33_ASAP7_75t_R      g285( .A (x51), .B (x179), .Y (n593) );
  AND2x2_ASAP7_75t_R        g286( .A (x51), .B (x179), .Y (n595) );
  NOR2xp33_ASAP7_75t_R      g287( .A (n593), .B (n595), .Y (n596) );
  XOR2xp5_ASAP7_75t_R       g288( .A (n592), .B (n596), .Y (y51) );
  OR2x2_ASAP7_75t_R         g289( .A (x52), .B (x180), .Y (n599) );
  NAND2xp33_ASAP7_75t_R     g290( .A (x52), .B (x180), .Y (n600) );
  NAND2xp33_ASAP7_75t_R     g291( .A (n599), .B (n600), .Y (n602) );
  INVx1_ASAP7_75t_R         g292( .A (n593), .Y (n594) );
  AOI21xp33_ASAP7_75t_R     g293( .A1 (n592), .B (n595), .A2 (n594), .Y (n598) );
  XOR2xp5_ASAP7_75t_R       g294( .A (n602), .B (n598), .Y (y52) );
  XNOR2xp5_ASAP7_75t_R      g295( .A (x53), .B (x181), .Y (n605) );
  INVx1_ASAP7_75t_R         g296( .A (n600), .Y (n601) );
  A2O1A1O1Ixp25_ASAP7_75t_R g297( .A1 (n592), .B (n595), .D (n601), .A2 (n594), .C (n599), .Y (n604) );
  XOR2xp5_ASAP7_75t_R       g298( .A (n605), .B (n604), .Y (y53) );
  INVx1_ASAP7_75t_R         g299( .A (x53), .Y (n274) );
  INVx1_ASAP7_75t_R         g300( .A (x181), .Y (n315) );
  MAJIxp5_ASAP7_75t_R       g301( .A (n274), .B (n315), .C (n604), .Y (n607) );
  NOR2xp33_ASAP7_75t_R      g302( .A (x54), .B (x182), .Y (n608) );
  AND2x2_ASAP7_75t_R        g303( .A (x54), .B (x182), .Y (n610) );
  NOR2xp33_ASAP7_75t_R      g304( .A (n608), .B (n610), .Y (n611) );
  XOR2xp5_ASAP7_75t_R       g305( .A (n607), .B (n611), .Y (y54) );
  OR2x2_ASAP7_75t_R         g306( .A (x55), .B (x183), .Y (n614) );
  NAND2xp33_ASAP7_75t_R     g307( .A (x55), .B (x183), .Y (n615) );
  NAND2xp33_ASAP7_75t_R     g308( .A (n614), .B (n615), .Y (n617) );
  INVx1_ASAP7_75t_R         g309( .A (n608), .Y (n609) );
  AOI21xp33_ASAP7_75t_R     g310( .A1 (n607), .B (n610), .A2 (n609), .Y (n613) );
  XOR2xp5_ASAP7_75t_R       g311( .A (n617), .B (n613), .Y (y55) );
  XNOR2xp5_ASAP7_75t_R      g312( .A (x56), .B (x184), .Y (n620) );
  INVx1_ASAP7_75t_R         g313( .A (n615), .Y (n616) );
  A2O1A1O1Ixp25_ASAP7_75t_R g314( .A1 (n607), .B (n610), .D (n616), .A2 (n609), .C (n614), .Y (n619) );
  XOR2xp5_ASAP7_75t_R       g315( .A (n620), .B (n619), .Y (y56) );
  INVx1_ASAP7_75t_R         g316( .A (x56), .Y (n275) );
  INVx1_ASAP7_75t_R         g317( .A (x184), .Y (n316) );
  MAJIxp5_ASAP7_75t_R       g318( .A (n275), .B (n316), .C (n619), .Y (n622) );
  NOR2xp33_ASAP7_75t_R      g319( .A (x57), .B (x185), .Y (n623) );
  AND2x2_ASAP7_75t_R        g320( .A (x57), .B (x185), .Y (n625) );
  NOR2xp33_ASAP7_75t_R      g321( .A (n623), .B (n625), .Y (n626) );
  XOR2xp5_ASAP7_75t_R       g322( .A (n622), .B (n626), .Y (y57) );
  OR2x2_ASAP7_75t_R         g323( .A (x58), .B (x186), .Y (n629) );
  NAND2xp33_ASAP7_75t_R     g324( .A (x58), .B (x186), .Y (n630) );
  NAND2xp33_ASAP7_75t_R     g325( .A (n629), .B (n630), .Y (n632) );
  INVx1_ASAP7_75t_R         g326( .A (n623), .Y (n624) );
  AOI21xp33_ASAP7_75t_R     g327( .A1 (n622), .B (n625), .A2 (n624), .Y (n628) );
  XOR2xp5_ASAP7_75t_R       g328( .A (n632), .B (n628), .Y (y58) );
  XNOR2xp5_ASAP7_75t_R      g329( .A (x59), .B (x187), .Y (n635) );
  INVx1_ASAP7_75t_R         g330( .A (n630), .Y (n631) );
  A2O1A1O1Ixp25_ASAP7_75t_R g331( .A1 (n622), .B (n625), .D (n631), .A2 (n624), .C (n629), .Y (n634) );
  XOR2xp5_ASAP7_75t_R       g332( .A (n635), .B (n634), .Y (y59) );
  INVx1_ASAP7_75t_R         g333( .A (x59), .Y (n276) );
  INVx1_ASAP7_75t_R         g334( .A (x187), .Y (n317) );
  MAJIxp5_ASAP7_75t_R       g335( .A (n276), .B (n317), .C (n634), .Y (n637) );
  NOR2xp33_ASAP7_75t_R      g336( .A (x60), .B (x188), .Y (n638) );
  AND2x2_ASAP7_75t_R        g337( .A (x60), .B (x188), .Y (n640) );
  NOR2xp33_ASAP7_75t_R      g338( .A (n638), .B (n640), .Y (n641) );
  XOR2xp5_ASAP7_75t_R       g339( .A (n637), .B (n641), .Y (y60) );
  OR2x2_ASAP7_75t_R         g340( .A (x61), .B (x189), .Y (n644) );
  NAND2xp33_ASAP7_75t_R     g341( .A (x61), .B (x189), .Y (n645) );
  NAND2xp33_ASAP7_75t_R     g342( .A (n644), .B (n645), .Y (n647) );
  INVx1_ASAP7_75t_R         g343( .A (n638), .Y (n639) );
  AOI21xp33_ASAP7_75t_R     g344( .A1 (n637), .B (n640), .A2 (n639), .Y (n643) );
  XOR2xp5_ASAP7_75t_R       g345( .A (n647), .B (n643), .Y (y61) );
  XNOR2xp5_ASAP7_75t_R      g346( .A (x62), .B (x190), .Y (n650) );
  INVx1_ASAP7_75t_R         g347( .A (n645), .Y (n646) );
  A2O1A1O1Ixp25_ASAP7_75t_R g348( .A1 (n637), .B (n640), .D (n646), .A2 (n639), .C (n644), .Y (n649) );
  XOR2xp5_ASAP7_75t_R       g349( .A (n650), .B (n649), .Y (y62) );
  INVx1_ASAP7_75t_R         g350( .A (x62), .Y (n277) );
  INVx1_ASAP7_75t_R         g351( .A (x190), .Y (n318) );
  MAJIxp5_ASAP7_75t_R       g352( .A (n277), .B (n318), .C (n649), .Y (n652) );
  NOR2xp33_ASAP7_75t_R      g353( .A (x63), .B (x191), .Y (n653) );
  AND2x2_ASAP7_75t_R        g354( .A (x63), .B (x191), .Y (n655) );
  NOR2xp33_ASAP7_75t_R      g355( .A (n653), .B (n655), .Y (n656) );
  XOR2xp5_ASAP7_75t_R       g356( .A (n652), .B (n656), .Y (y63) );
  OR2x2_ASAP7_75t_R         g357( .A (x64), .B (x192), .Y (n659) );
  NAND2xp33_ASAP7_75t_R     g358( .A (x64), .B (x192), .Y (n660) );
  NAND2xp33_ASAP7_75t_R     g359( .A (n659), .B (n660), .Y (n662) );
  INVx1_ASAP7_75t_R         g360( .A (n653), .Y (n654) );
  AOI21xp33_ASAP7_75t_R     g361( .A1 (n652), .B (n655), .A2 (n654), .Y (n658) );
  XOR2xp5_ASAP7_75t_R       g362( .A (n662), .B (n658), .Y (y64) );
  XNOR2xp5_ASAP7_75t_R      g363( .A (x65), .B (x193), .Y (n665) );
  INVx1_ASAP7_75t_R         g364( .A (n660), .Y (n661) );
  A2O1A1O1Ixp25_ASAP7_75t_R g365( .A1 (n652), .B (n655), .D (n661), .A2 (n654), .C (n659), .Y (n664) );
  XOR2xp5_ASAP7_75t_R       g366( .A (n665), .B (n664), .Y (y65) );
  INVx1_ASAP7_75t_R         g367( .A (x65), .Y (n278) );
  INVx1_ASAP7_75t_R         g368( .A (x193), .Y (n319) );
  MAJIxp5_ASAP7_75t_R       g369( .A (n278), .B (n319), .C (n664), .Y (n667) );
  NOR2xp33_ASAP7_75t_R      g370( .A (x66), .B (x194), .Y (n668) );
  AND2x2_ASAP7_75t_R        g371( .A (x66), .B (x194), .Y (n670) );
  NOR2xp33_ASAP7_75t_R      g372( .A (n668), .B (n670), .Y (n671) );
  XOR2xp5_ASAP7_75t_R       g373( .A (n667), .B (n671), .Y (y66) );
  OR2x2_ASAP7_75t_R         g374( .A (x67), .B (x195), .Y (n674) );
  NAND2xp33_ASAP7_75t_R     g375( .A (x67), .B (x195), .Y (n675) );
  NAND2xp33_ASAP7_75t_R     g376( .A (n674), .B (n675), .Y (n677) );
  INVx1_ASAP7_75t_R         g377( .A (n668), .Y (n669) );
  AOI21xp33_ASAP7_75t_R     g378( .A1 (n667), .B (n670), .A2 (n669), .Y (n673) );
  XOR2xp5_ASAP7_75t_R       g379( .A (n677), .B (n673), .Y (y67) );
  XNOR2xp5_ASAP7_75t_R      g380( .A (x68), .B (x196), .Y (n680) );
  INVx1_ASAP7_75t_R         g381( .A (n675), .Y (n676) );
  A2O1A1O1Ixp25_ASAP7_75t_R g382( .A1 (n667), .B (n670), .D (n676), .A2 (n669), .C (n674), .Y (n679) );
  XOR2xp5_ASAP7_75t_R       g383( .A (n680), .B (n679), .Y (y68) );
  INVx1_ASAP7_75t_R         g384( .A (x68), .Y (n279) );
  INVx1_ASAP7_75t_R         g385( .A (x196), .Y (n320) );
  MAJIxp5_ASAP7_75t_R       g386( .A (n279), .B (n320), .C (n679), .Y (n682) );
  NOR2xp33_ASAP7_75t_R      g387( .A (x69), .B (x197), .Y (n683) );
  AND2x2_ASAP7_75t_R        g388( .A (x69), .B (x197), .Y (n685) );
  NOR2xp33_ASAP7_75t_R      g389( .A (n683), .B (n685), .Y (n686) );
  XOR2xp5_ASAP7_75t_R       g390( .A (n682), .B (n686), .Y (y69) );
  OR2x2_ASAP7_75t_R         g391( .A (x70), .B (x198), .Y (n689) );
  NAND2xp33_ASAP7_75t_R     g392( .A (x70), .B (x198), .Y (n690) );
  NAND2xp33_ASAP7_75t_R     g393( .A (n689), .B (n690), .Y (n692) );
  INVx1_ASAP7_75t_R         g394( .A (n683), .Y (n684) );
  AOI21xp33_ASAP7_75t_R     g395( .A1 (n682), .B (n685), .A2 (n684), .Y (n688) );
  XOR2xp5_ASAP7_75t_R       g396( .A (n692), .B (n688), .Y (y70) );
  XNOR2xp5_ASAP7_75t_R      g397( .A (x71), .B (x199), .Y (n695) );
  INVx1_ASAP7_75t_R         g398( .A (n690), .Y (n691) );
  A2O1A1O1Ixp25_ASAP7_75t_R g399( .A1 (n682), .B (n685), .D (n691), .A2 (n684), .C (n689), .Y (n694) );
  XOR2xp5_ASAP7_75t_R       g400( .A (n695), .B (n694), .Y (y71) );
  INVx1_ASAP7_75t_R         g401( .A (x71), .Y (n280) );
  INVx1_ASAP7_75t_R         g402( .A (x199), .Y (n321) );
  MAJIxp5_ASAP7_75t_R       g403( .A (n280), .B (n321), .C (n694), .Y (n697) );
  NOR2xp33_ASAP7_75t_R      g404( .A (x72), .B (x200), .Y (n698) );
  AND2x2_ASAP7_75t_R        g405( .A (x72), .B (x200), .Y (n700) );
  NOR2xp33_ASAP7_75t_R      g406( .A (n698), .B (n700), .Y (n701) );
  XOR2xp5_ASAP7_75t_R       g407( .A (n697), .B (n701), .Y (y72) );
  OR2x2_ASAP7_75t_R         g408( .A (x73), .B (x201), .Y (n704) );
  NAND2xp33_ASAP7_75t_R     g409( .A (x73), .B (x201), .Y (n705) );
  NAND2xp33_ASAP7_75t_R     g410( .A (n704), .B (n705), .Y (n707) );
  INVx1_ASAP7_75t_R         g411( .A (n698), .Y (n699) );
  AOI21xp33_ASAP7_75t_R     g412( .A1 (n697), .B (n700), .A2 (n699), .Y (n703) );
  XOR2xp5_ASAP7_75t_R       g413( .A (n707), .B (n703), .Y (y73) );
  XNOR2xp5_ASAP7_75t_R      g414( .A (x74), .B (x202), .Y (n710) );
  INVx1_ASAP7_75t_R         g415( .A (n705), .Y (n706) );
  A2O1A1O1Ixp25_ASAP7_75t_R g416( .A1 (n697), .B (n700), .D (n706), .A2 (n699), .C (n704), .Y (n709) );
  XOR2xp5_ASAP7_75t_R       g417( .A (n710), .B (n709), .Y (y74) );
  INVx1_ASAP7_75t_R         g418( .A (x74), .Y (n281) );
  INVx1_ASAP7_75t_R         g419( .A (x202), .Y (n322) );
  MAJIxp5_ASAP7_75t_R       g420( .A (n281), .B (n322), .C (n709), .Y (n712) );
  NOR2xp33_ASAP7_75t_R      g421( .A (x75), .B (x203), .Y (n713) );
  AND2x2_ASAP7_75t_R        g422( .A (x75), .B (x203), .Y (n715) );
  NOR2xp33_ASAP7_75t_R      g423( .A (n713), .B (n715), .Y (n716) );
  XOR2xp5_ASAP7_75t_R       g424( .A (n712), .B (n716), .Y (y75) );
  OR2x2_ASAP7_75t_R         g425( .A (x76), .B (x204), .Y (n719) );
  NAND2xp33_ASAP7_75t_R     g426( .A (x76), .B (x204), .Y (n720) );
  NAND2xp33_ASAP7_75t_R     g427( .A (n719), .B (n720), .Y (n722) );
  INVx1_ASAP7_75t_R         g428( .A (n713), .Y (n714) );
  AOI21xp33_ASAP7_75t_R     g429( .A1 (n712), .B (n715), .A2 (n714), .Y (n718) );
  XOR2xp5_ASAP7_75t_R       g430( .A (n722), .B (n718), .Y (y76) );
  XNOR2xp5_ASAP7_75t_R      g431( .A (x77), .B (x205), .Y (n725) );
  INVx1_ASAP7_75t_R         g432( .A (n720), .Y (n721) );
  A2O1A1O1Ixp25_ASAP7_75t_R g433( .A1 (n712), .B (n715), .D (n721), .A2 (n714), .C (n719), .Y (n724) );
  XOR2xp5_ASAP7_75t_R       g434( .A (n725), .B (n724), .Y (y77) );
  INVx1_ASAP7_75t_R         g435( .A (x77), .Y (n282) );
  INVx1_ASAP7_75t_R         g436( .A (x205), .Y (n323) );
  MAJIxp5_ASAP7_75t_R       g437( .A (n282), .B (n323), .C (n724), .Y (n727) );
  NOR2xp33_ASAP7_75t_R      g438( .A (x78), .B (x206), .Y (n728) );
  AND2x2_ASAP7_75t_R        g439( .A (x78), .B (x206), .Y (n730) );
  NOR2xp33_ASAP7_75t_R      g440( .A (n728), .B (n730), .Y (n731) );
  XOR2xp5_ASAP7_75t_R       g441( .A (n727), .B (n731), .Y (y78) );
  OR2x2_ASAP7_75t_R         g442( .A (x79), .B (x207), .Y (n734) );
  NAND2xp33_ASAP7_75t_R     g443( .A (x79), .B (x207), .Y (n735) );
  NAND2xp33_ASAP7_75t_R     g444( .A (n734), .B (n735), .Y (n737) );
  INVx1_ASAP7_75t_R         g445( .A (n728), .Y (n729) );
  AOI21xp33_ASAP7_75t_R     g446( .A1 (n727), .B (n730), .A2 (n729), .Y (n733) );
  XOR2xp5_ASAP7_75t_R       g447( .A (n737), .B (n733), .Y (y79) );
  XNOR2xp5_ASAP7_75t_R      g448( .A (x80), .B (x208), .Y (n740) );
  INVx1_ASAP7_75t_R         g449( .A (n735), .Y (n736) );
  A2O1A1O1Ixp25_ASAP7_75t_R g450( .A1 (n727), .B (n730), .D (n736), .A2 (n729), .C (n734), .Y (n739) );
  XOR2xp5_ASAP7_75t_R       g451( .A (n740), .B (n739), .Y (y80) );
  INVx1_ASAP7_75t_R         g452( .A (x80), .Y (n283) );
  INVx1_ASAP7_75t_R         g453( .A (x208), .Y (n324) );
  MAJIxp5_ASAP7_75t_R       g454( .A (n283), .B (n324), .C (n739), .Y (n742) );
  NOR2xp33_ASAP7_75t_R      g455( .A (x81), .B (x209), .Y (n743) );
  AND2x2_ASAP7_75t_R        g456( .A (x81), .B (x209), .Y (n745) );
  NOR2xp33_ASAP7_75t_R      g457( .A (n743), .B (n745), .Y (n746) );
  XOR2xp5_ASAP7_75t_R       g458( .A (n742), .B (n746), .Y (y81) );
  OR2x2_ASAP7_75t_R         g459( .A (x82), .B (x210), .Y (n749) );
  NAND2xp33_ASAP7_75t_R     g460( .A (x82), .B (x210), .Y (n750) );
  NAND2xp33_ASAP7_75t_R     g461( .A (n749), .B (n750), .Y (n752) );
  INVx1_ASAP7_75t_R         g462( .A (n743), .Y (n744) );
  AOI21xp33_ASAP7_75t_R     g463( .A1 (n742), .B (n745), .A2 (n744), .Y (n748) );
  XOR2xp5_ASAP7_75t_R       g464( .A (n752), .B (n748), .Y (y82) );
  XNOR2xp5_ASAP7_75t_R      g465( .A (x83), .B (x211), .Y (n755) );
  INVx1_ASAP7_75t_R         g466( .A (n750), .Y (n751) );
  A2O1A1O1Ixp25_ASAP7_75t_R g467( .A1 (n742), .B (n745), .D (n751), .A2 (n744), .C (n749), .Y (n754) );
  XOR2xp5_ASAP7_75t_R       g468( .A (n755), .B (n754), .Y (y83) );
  INVx1_ASAP7_75t_R         g469( .A (x83), .Y (n284) );
  INVx1_ASAP7_75t_R         g470( .A (x211), .Y (n325) );
  MAJIxp5_ASAP7_75t_R       g471( .A (n284), .B (n325), .C (n754), .Y (n757) );
  NOR2xp33_ASAP7_75t_R      g472( .A (x84), .B (x212), .Y (n758) );
  AND2x2_ASAP7_75t_R        g473( .A (x84), .B (x212), .Y (n760) );
  NOR2xp33_ASAP7_75t_R      g474( .A (n758), .B (n760), .Y (n761) );
  XOR2xp5_ASAP7_75t_R       g475( .A (n757), .B (n761), .Y (y84) );
  OR2x2_ASAP7_75t_R         g476( .A (x85), .B (x213), .Y (n764) );
  NAND2xp33_ASAP7_75t_R     g477( .A (x85), .B (x213), .Y (n765) );
  NAND2xp33_ASAP7_75t_R     g478( .A (n764), .B (n765), .Y (n767) );
  INVx1_ASAP7_75t_R         g479( .A (n758), .Y (n759) );
  AOI21xp33_ASAP7_75t_R     g480( .A1 (n757), .B (n760), .A2 (n759), .Y (n763) );
  XOR2xp5_ASAP7_75t_R       g481( .A (n767), .B (n763), .Y (y85) );
  XNOR2xp5_ASAP7_75t_R      g482( .A (x86), .B (x214), .Y (n770) );
  INVx1_ASAP7_75t_R         g483( .A (n765), .Y (n766) );
  A2O1A1O1Ixp25_ASAP7_75t_R g484( .A1 (n757), .B (n760), .D (n766), .A2 (n759), .C (n764), .Y (n769) );
  XOR2xp5_ASAP7_75t_R       g485( .A (n770), .B (n769), .Y (y86) );
  INVx1_ASAP7_75t_R         g486( .A (x86), .Y (n285) );
  INVx1_ASAP7_75t_R         g487( .A (x214), .Y (n326) );
  MAJIxp5_ASAP7_75t_R       g488( .A (n285), .B (n326), .C (n769), .Y (n772) );
  NOR2xp33_ASAP7_75t_R      g489( .A (x87), .B (x215), .Y (n773) );
  AND2x2_ASAP7_75t_R        g490( .A (x87), .B (x215), .Y (n775) );
  NOR2xp33_ASAP7_75t_R      g491( .A (n773), .B (n775), .Y (n776) );
  XOR2xp5_ASAP7_75t_R       g492( .A (n772), .B (n776), .Y (y87) );
  OR2x2_ASAP7_75t_R         g493( .A (x88), .B (x216), .Y (n779) );
  NAND2xp33_ASAP7_75t_R     g494( .A (x88), .B (x216), .Y (n780) );
  NAND2xp33_ASAP7_75t_R     g495( .A (n779), .B (n780), .Y (n782) );
  INVx1_ASAP7_75t_R         g496( .A (n773), .Y (n774) );
  AOI21xp33_ASAP7_75t_R     g497( .A1 (n772), .B (n775), .A2 (n774), .Y (n778) );
  XOR2xp5_ASAP7_75t_R       g498( .A (n782), .B (n778), .Y (y88) );
  XNOR2xp5_ASAP7_75t_R      g499( .A (x89), .B (x217), .Y (n785) );
  INVx1_ASAP7_75t_R         g500( .A (n780), .Y (n781) );
  A2O1A1O1Ixp25_ASAP7_75t_R g501( .A1 (n772), .B (n775), .D (n781), .A2 (n774), .C (n779), .Y (n784) );
  XOR2xp5_ASAP7_75t_R       g502( .A (n785), .B (n784), .Y (y89) );
  INVx1_ASAP7_75t_R         g503( .A (x89), .Y (n286) );
  INVx1_ASAP7_75t_R         g504( .A (x217), .Y (n327) );
  MAJIxp5_ASAP7_75t_R       g505( .A (n286), .B (n327), .C (n784), .Y (n787) );
  NOR2xp33_ASAP7_75t_R      g506( .A (x90), .B (x218), .Y (n788) );
  AND2x2_ASAP7_75t_R        g507( .A (x90), .B (x218), .Y (n790) );
  NOR2xp33_ASAP7_75t_R      g508( .A (n788), .B (n790), .Y (n791) );
  XOR2xp5_ASAP7_75t_R       g509( .A (n787), .B (n791), .Y (y90) );
  OR2x2_ASAP7_75t_R         g510( .A (x91), .B (x219), .Y (n794) );
  NAND2xp33_ASAP7_75t_R     g511( .A (x91), .B (x219), .Y (n795) );
  NAND2xp33_ASAP7_75t_R     g512( .A (n794), .B (n795), .Y (n797) );
  INVx1_ASAP7_75t_R         g513( .A (n788), .Y (n789) );
  AOI21xp33_ASAP7_75t_R     g514( .A1 (n787), .B (n790), .A2 (n789), .Y (n793) );
  XOR2xp5_ASAP7_75t_R       g515( .A (n797), .B (n793), .Y (y91) );
  XNOR2xp5_ASAP7_75t_R      g516( .A (x92), .B (x220), .Y (n800) );
  INVx1_ASAP7_75t_R         g517( .A (n795), .Y (n796) );
  A2O1A1O1Ixp25_ASAP7_75t_R g518( .A1 (n787), .B (n790), .D (n796), .A2 (n789), .C (n794), .Y (n799) );
  XOR2xp5_ASAP7_75t_R       g519( .A (n800), .B (n799), .Y (y92) );
  INVx1_ASAP7_75t_R         g520( .A (x92), .Y (n287) );
  INVx1_ASAP7_75t_R         g521( .A (x220), .Y (n328) );
  MAJIxp5_ASAP7_75t_R       g522( .A (n287), .B (n328), .C (n799), .Y (n802) );
  NOR2xp33_ASAP7_75t_R      g523( .A (x93), .B (x221), .Y (n803) );
  AND2x2_ASAP7_75t_R        g524( .A (x93), .B (x221), .Y (n805) );
  NOR2xp33_ASAP7_75t_R      g525( .A (n803), .B (n805), .Y (n806) );
  XOR2xp5_ASAP7_75t_R       g526( .A (n802), .B (n806), .Y (y93) );
  OR2x2_ASAP7_75t_R         g527( .A (x94), .B (x222), .Y (n809) );
  NAND2xp33_ASAP7_75t_R     g528( .A (x94), .B (x222), .Y (n810) );
  NAND2xp33_ASAP7_75t_R     g529( .A (n809), .B (n810), .Y (n812) );
  INVx1_ASAP7_75t_R         g530( .A (n803), .Y (n804) );
  AOI21xp33_ASAP7_75t_R     g531( .A1 (n802), .B (n805), .A2 (n804), .Y (n808) );
  XOR2xp5_ASAP7_75t_R       g532( .A (n812), .B (n808), .Y (y94) );
  XNOR2xp5_ASAP7_75t_R      g533( .A (x95), .B (x223), .Y (n815) );
  INVx1_ASAP7_75t_R         g534( .A (n810), .Y (n811) );
  A2O1A1O1Ixp25_ASAP7_75t_R g535( .A1 (n802), .B (n805), .D (n811), .A2 (n804), .C (n809), .Y (n814) );
  XOR2xp5_ASAP7_75t_R       g536( .A (n815), .B (n814), .Y (y95) );
  INVx1_ASAP7_75t_R         g537( .A (x95), .Y (n288) );
  INVx1_ASAP7_75t_R         g538( .A (x223), .Y (n329) );
  MAJIxp5_ASAP7_75t_R       g539( .A (n288), .B (n329), .C (n814), .Y (n817) );
  NOR2xp33_ASAP7_75t_R      g540( .A (x96), .B (x224), .Y (n818) );
  AND2x2_ASAP7_75t_R        g541( .A (x96), .B (x224), .Y (n820) );
  NOR2xp33_ASAP7_75t_R      g542( .A (n818), .B (n820), .Y (n821) );
  XOR2xp5_ASAP7_75t_R       g543( .A (n817), .B (n821), .Y (y96) );
  OR2x2_ASAP7_75t_R         g544( .A (x97), .B (x225), .Y (n824) );
  NAND2xp33_ASAP7_75t_R     g545( .A (x97), .B (x225), .Y (n825) );
  NAND2xp33_ASAP7_75t_R     g546( .A (n824), .B (n825), .Y (n827) );
  INVx1_ASAP7_75t_R         g547( .A (n818), .Y (n819) );
  AOI21xp33_ASAP7_75t_R     g548( .A1 (n817), .B (n820), .A2 (n819), .Y (n823) );
  XOR2xp5_ASAP7_75t_R       g549( .A (n827), .B (n823), .Y (y97) );
  XNOR2xp5_ASAP7_75t_R      g550( .A (x98), .B (x226), .Y (n830) );
  INVx1_ASAP7_75t_R         g551( .A (n825), .Y (n826) );
  A2O1A1O1Ixp25_ASAP7_75t_R g552( .A1 (n817), .B (n820), .D (n826), .A2 (n819), .C (n824), .Y (n829) );
  XOR2xp5_ASAP7_75t_R       g553( .A (n830), .B (n829), .Y (y98) );
  INVx1_ASAP7_75t_R         g554( .A (x98), .Y (n289) );
  INVx1_ASAP7_75t_R         g555( .A (x226), .Y (n330) );
  MAJIxp5_ASAP7_75t_R       g556( .A (n289), .B (n330), .C (n829), .Y (n832) );
  NOR2xp33_ASAP7_75t_R      g557( .A (x99), .B (x227), .Y (n833) );
  AND2x2_ASAP7_75t_R        g558( .A (x99), .B (x227), .Y (n835) );
  NOR2xp33_ASAP7_75t_R      g559( .A (n833), .B (n835), .Y (n836) );
  XOR2xp5_ASAP7_75t_R       g560( .A (n832), .B (n836), .Y (y99) );
  OR2x2_ASAP7_75t_R         g561( .A (x100), .B (x228), .Y (n839) );
  NAND2xp33_ASAP7_75t_R     g562( .A (x100), .B (x228), .Y (n840) );
  NAND2xp33_ASAP7_75t_R     g563( .A (n839), .B (n840), .Y (n842) );
  INVx1_ASAP7_75t_R         g564( .A (n833), .Y (n834) );
  AOI21xp33_ASAP7_75t_R     g565( .A1 (n832), .B (n835), .A2 (n834), .Y (n838) );
  XOR2xp5_ASAP7_75t_R       g566( .A (n842), .B (n838), .Y (y100) );
  XNOR2xp5_ASAP7_75t_R      g567( .A (x101), .B (x229), .Y (n845) );
  INVx1_ASAP7_75t_R         g568( .A (n840), .Y (n841) );
  A2O1A1O1Ixp25_ASAP7_75t_R g569( .A1 (n832), .B (n835), .D (n841), .A2 (n834), .C (n839), .Y (n844) );
  XOR2xp5_ASAP7_75t_R       g570( .A (n845), .B (n844), .Y (y101) );
  INVx1_ASAP7_75t_R         g571( .A (x101), .Y (n290) );
  INVx1_ASAP7_75t_R         g572( .A (x229), .Y (n331) );
  MAJIxp5_ASAP7_75t_R       g573( .A (n290), .B (n331), .C (n844), .Y (n847) );
  NOR2xp33_ASAP7_75t_R      g574( .A (x102), .B (x230), .Y (n848) );
  AND2x2_ASAP7_75t_R        g575( .A (x102), .B (x230), .Y (n850) );
  NOR2xp33_ASAP7_75t_R      g576( .A (n848), .B (n850), .Y (n851) );
  XOR2xp5_ASAP7_75t_R       g577( .A (n847), .B (n851), .Y (y102) );
  OR2x2_ASAP7_75t_R         g578( .A (x103), .B (x231), .Y (n854) );
  NAND2xp33_ASAP7_75t_R     g579( .A (x103), .B (x231), .Y (n855) );
  NAND2xp33_ASAP7_75t_R     g580( .A (n854), .B (n855), .Y (n857) );
  INVx1_ASAP7_75t_R         g581( .A (n848), .Y (n849) );
  AOI21xp33_ASAP7_75t_R     g582( .A1 (n847), .B (n850), .A2 (n849), .Y (n853) );
  XOR2xp5_ASAP7_75t_R       g583( .A (n857), .B (n853), .Y (y103) );
  XNOR2xp5_ASAP7_75t_R      g584( .A (x104), .B (x232), .Y (n860) );
  INVx1_ASAP7_75t_R         g585( .A (n855), .Y (n856) );
  A2O1A1O1Ixp25_ASAP7_75t_R g586( .A1 (n847), .B (n850), .D (n856), .A2 (n849), .C (n854), .Y (n859) );
  XOR2xp5_ASAP7_75t_R       g587( .A (n860), .B (n859), .Y (y104) );
  INVx1_ASAP7_75t_R         g588( .A (x104), .Y (n291) );
  INVx1_ASAP7_75t_R         g589( .A (x232), .Y (n332) );
  MAJIxp5_ASAP7_75t_R       g590( .A (n291), .B (n332), .C (n859), .Y (n862) );
  NOR2xp33_ASAP7_75t_R      g591( .A (x105), .B (x233), .Y (n863) );
  AND2x2_ASAP7_75t_R        g592( .A (x105), .B (x233), .Y (n865) );
  NOR2xp33_ASAP7_75t_R      g593( .A (n863), .B (n865), .Y (n866) );
  XOR2xp5_ASAP7_75t_R       g594( .A (n862), .B (n866), .Y (y105) );
  OR2x2_ASAP7_75t_R         g595( .A (x106), .B (x234), .Y (n869) );
  NAND2xp33_ASAP7_75t_R     g596( .A (x106), .B (x234), .Y (n870) );
  NAND2xp33_ASAP7_75t_R     g597( .A (n869), .B (n870), .Y (n872) );
  INVx1_ASAP7_75t_R         g598( .A (n863), .Y (n864) );
  AOI21xp33_ASAP7_75t_R     g599( .A1 (n862), .B (n865), .A2 (n864), .Y (n868) );
  XOR2xp5_ASAP7_75t_R       g600( .A (n872), .B (n868), .Y (y106) );
  XNOR2xp5_ASAP7_75t_R      g601( .A (x107), .B (x235), .Y (n875) );
  INVx1_ASAP7_75t_R         g602( .A (n870), .Y (n871) );
  A2O1A1O1Ixp25_ASAP7_75t_R g603( .A1 (n862), .B (n865), .D (n871), .A2 (n864), .C (n869), .Y (n874) );
  XOR2xp5_ASAP7_75t_R       g604( .A (n875), .B (n874), .Y (y107) );
  INVx1_ASAP7_75t_R         g605( .A (x107), .Y (n292) );
  INVx1_ASAP7_75t_R         g606( .A (x235), .Y (n333) );
  MAJIxp5_ASAP7_75t_R       g607( .A (n292), .B (n333), .C (n874), .Y (n877) );
  NOR2xp33_ASAP7_75t_R      g608( .A (x108), .B (x236), .Y (n878) );
  AND2x2_ASAP7_75t_R        g609( .A (x108), .B (x236), .Y (n880) );
  NOR2xp33_ASAP7_75t_R      g610( .A (n878), .B (n880), .Y (n881) );
  XOR2xp5_ASAP7_75t_R       g611( .A (n877), .B (n881), .Y (y108) );
  OR2x2_ASAP7_75t_R         g612( .A (x109), .B (x237), .Y (n884) );
  NAND2xp33_ASAP7_75t_R     g613( .A (x109), .B (x237), .Y (n885) );
  NAND2xp33_ASAP7_75t_R     g614( .A (n884), .B (n885), .Y (n887) );
  INVx1_ASAP7_75t_R         g615( .A (n878), .Y (n879) );
  AOI21xp33_ASAP7_75t_R     g616( .A1 (n877), .B (n880), .A2 (n879), .Y (n883) );
  XOR2xp5_ASAP7_75t_R       g617( .A (n887), .B (n883), .Y (y109) );
  XNOR2xp5_ASAP7_75t_R      g618( .A (x110), .B (x238), .Y (n890) );
  INVx1_ASAP7_75t_R         g619( .A (n885), .Y (n886) );
  A2O1A1O1Ixp25_ASAP7_75t_R g620( .A1 (n877), .B (n880), .D (n886), .A2 (n879), .C (n884), .Y (n889) );
  XOR2xp5_ASAP7_75t_R       g621( .A (n890), .B (n889), .Y (y110) );
  INVx1_ASAP7_75t_R         g622( .A (x110), .Y (n293) );
  INVx1_ASAP7_75t_R         g623( .A (x238), .Y (n334) );
  MAJIxp5_ASAP7_75t_R       g624( .A (n293), .B (n334), .C (n889), .Y (n892) );
  NOR2xp33_ASAP7_75t_R      g625( .A (x111), .B (x239), .Y (n893) );
  AND2x2_ASAP7_75t_R        g626( .A (x111), .B (x239), .Y (n895) );
  NOR2xp33_ASAP7_75t_R      g627( .A (n893), .B (n895), .Y (n896) );
  XOR2xp5_ASAP7_75t_R       g628( .A (n892), .B (n896), .Y (y111) );
  OR2x2_ASAP7_75t_R         g629( .A (x112), .B (x240), .Y (n899) );
  NAND2xp33_ASAP7_75t_R     g630( .A (x112), .B (x240), .Y (n900) );
  NAND2xp33_ASAP7_75t_R     g631( .A (n899), .B (n900), .Y (n902) );
  INVx1_ASAP7_75t_R         g632( .A (n893), .Y (n894) );
  AOI21xp33_ASAP7_75t_R     g633( .A1 (n892), .B (n895), .A2 (n894), .Y (n898) );
  XOR2xp5_ASAP7_75t_R       g634( .A (n902), .B (n898), .Y (y112) );
  XNOR2xp5_ASAP7_75t_R      g635( .A (x113), .B (x241), .Y (n905) );
  INVx1_ASAP7_75t_R         g636( .A (n900), .Y (n901) );
  A2O1A1O1Ixp25_ASAP7_75t_R g637( .A1 (n892), .B (n895), .D (n901), .A2 (n894), .C (n899), .Y (n904) );
  XOR2xp5_ASAP7_75t_R       g638( .A (n905), .B (n904), .Y (y113) );
  INVx1_ASAP7_75t_R         g639( .A (x113), .Y (n294) );
  INVx1_ASAP7_75t_R         g640( .A (x241), .Y (n335) );
  MAJIxp5_ASAP7_75t_R       g641( .A (n294), .B (n335), .C (n904), .Y (n907) );
  NOR2xp33_ASAP7_75t_R      g642( .A (x114), .B (x242), .Y (n908) );
  AND2x2_ASAP7_75t_R        g643( .A (x114), .B (x242), .Y (n910) );
  NOR2xp33_ASAP7_75t_R      g644( .A (n908), .B (n910), .Y (n911) );
  XOR2xp5_ASAP7_75t_R       g645( .A (n907), .B (n911), .Y (y114) );
  OR2x2_ASAP7_75t_R         g646( .A (x115), .B (x243), .Y (n914) );
  NAND2xp33_ASAP7_75t_R     g647( .A (x115), .B (x243), .Y (n915) );
  NAND2xp33_ASAP7_75t_R     g648( .A (n914), .B (n915), .Y (n917) );
  INVx1_ASAP7_75t_R         g649( .A (n908), .Y (n909) );
  AOI21xp33_ASAP7_75t_R     g650( .A1 (n907), .B (n910), .A2 (n909), .Y (n913) );
  XOR2xp5_ASAP7_75t_R       g651( .A (n917), .B (n913), .Y (y115) );
  XNOR2xp5_ASAP7_75t_R      g652( .A (x116), .B (x244), .Y (n920) );
  INVx1_ASAP7_75t_R         g653( .A (n915), .Y (n916) );
  A2O1A1O1Ixp25_ASAP7_75t_R g654( .A1 (n907), .B (n910), .D (n916), .A2 (n909), .C (n914), .Y (n919) );
  XOR2xp5_ASAP7_75t_R       g655( .A (n920), .B (n919), .Y (y116) );
  INVx1_ASAP7_75t_R         g656( .A (x116), .Y (n295) );
  INVx1_ASAP7_75t_R         g657( .A (x244), .Y (n336) );
  MAJIxp5_ASAP7_75t_R       g658( .A (n295), .B (n336), .C (n919), .Y (n922) );
  NOR2xp33_ASAP7_75t_R      g659( .A (x117), .B (x245), .Y (n923) );
  AND2x2_ASAP7_75t_R        g660( .A (x117), .B (x245), .Y (n925) );
  NOR2xp33_ASAP7_75t_R      g661( .A (n923), .B (n925), .Y (n926) );
  XOR2xp5_ASAP7_75t_R       g662( .A (n922), .B (n926), .Y (y117) );
  OR2x2_ASAP7_75t_R         g663( .A (x118), .B (x246), .Y (n929) );
  NAND2xp33_ASAP7_75t_R     g664( .A (x118), .B (x246), .Y (n930) );
  NAND2xp33_ASAP7_75t_R     g665( .A (n929), .B (n930), .Y (n932) );
  INVx1_ASAP7_75t_R         g666( .A (n923), .Y (n924) );
  AOI21xp33_ASAP7_75t_R     g667( .A1 (n922), .B (n925), .A2 (n924), .Y (n928) );
  XOR2xp5_ASAP7_75t_R       g668( .A (n932), .B (n928), .Y (y118) );
  XNOR2xp5_ASAP7_75t_R      g669( .A (x119), .B (x247), .Y (n935) );
  INVx1_ASAP7_75t_R         g670( .A (n930), .Y (n931) );
  A2O1A1O1Ixp25_ASAP7_75t_R g671( .A1 (n922), .B (n925), .D (n931), .A2 (n924), .C (n929), .Y (n934) );
  XOR2xp5_ASAP7_75t_R       g672( .A (n935), .B (n934), .Y (y119) );
  INVx1_ASAP7_75t_R         g673( .A (x119), .Y (n296) );
  INVx1_ASAP7_75t_R         g674( .A (x247), .Y (n337) );
  MAJIxp5_ASAP7_75t_R       g675( .A (n296), .B (n337), .C (n934), .Y (n937) );
  NOR2xp33_ASAP7_75t_R      g676( .A (x120), .B (x248), .Y (n938) );
  AND2x2_ASAP7_75t_R        g677( .A (x120), .B (x248), .Y (n940) );
  NOR2xp33_ASAP7_75t_R      g678( .A (n938), .B (n940), .Y (n941) );
  XOR2xp5_ASAP7_75t_R       g679( .A (n937), .B (n941), .Y (y120) );
  OR2x2_ASAP7_75t_R         g680( .A (x121), .B (x249), .Y (n944) );
  NAND2xp33_ASAP7_75t_R     g681( .A (x121), .B (x249), .Y (n945) );
  NAND2xp33_ASAP7_75t_R     g682( .A (n944), .B (n945), .Y (n947) );
  INVx1_ASAP7_75t_R         g683( .A (n938), .Y (n939) );
  AOI21xp33_ASAP7_75t_R     g684( .A1 (n937), .B (n940), .A2 (n939), .Y (n943) );
  XOR2xp5_ASAP7_75t_R       g685( .A (n947), .B (n943), .Y (y121) );
  XNOR2xp5_ASAP7_75t_R      g686( .A (x122), .B (x250), .Y (n950) );
  INVx1_ASAP7_75t_R         g687( .A (n945), .Y (n946) );
  A2O1A1O1Ixp25_ASAP7_75t_R g688( .A1 (n937), .B (n940), .D (n946), .A2 (n939), .C (n944), .Y (n949) );
  XOR2xp5_ASAP7_75t_R       g689( .A (n950), .B (n949), .Y (y122) );
  INVx1_ASAP7_75t_R         g690( .A (x122), .Y (n297) );
  INVx1_ASAP7_75t_R         g691( .A (x250), .Y (n338) );
  MAJIxp5_ASAP7_75t_R       g692( .A (n297), .B (n338), .C (n949), .Y (n952) );
  NOR2xp33_ASAP7_75t_R      g693( .A (x123), .B (x251), .Y (n953) );
  AND2x2_ASAP7_75t_R        g694( .A (x123), .B (x251), .Y (n955) );
  NOR2xp33_ASAP7_75t_R      g695( .A (n953), .B (n955), .Y (n956) );
  XOR2xp5_ASAP7_75t_R       g696( .A (n952), .B (n956), .Y (y123) );
  OR2x2_ASAP7_75t_R         g697( .A (x124), .B (x252), .Y (n959) );
  NAND2xp33_ASAP7_75t_R     g698( .A (x124), .B (x252), .Y (n960) );
  NAND2xp33_ASAP7_75t_R     g699( .A (n959), .B (n960), .Y (n962) );
  INVx1_ASAP7_75t_R         g700( .A (n953), .Y (n954) );
  AOI21xp33_ASAP7_75t_R     g701( .A1 (n952), .B (n955), .A2 (n954), .Y (n958) );
  XOR2xp5_ASAP7_75t_R       g702( .A (n962), .B (n958), .Y (y124) );
  XNOR2xp5_ASAP7_75t_R      g703( .A (x125), .B (x253), .Y (n965) );
  INVx1_ASAP7_75t_R         g704( .A (n960), .Y (n961) );
  A2O1A1O1Ixp25_ASAP7_75t_R g705( .A1 (n952), .B (n955), .D (n961), .A2 (n954), .C (n959), .Y (n964) );
  XOR2xp5_ASAP7_75t_R       g706( .A (n965), .B (n964), .Y (y125) );
  INVx1_ASAP7_75t_R         g707( .A (x125), .Y (n298) );
  INVx1_ASAP7_75t_R         g708( .A (x253), .Y (n339) );
  MAJIxp5_ASAP7_75t_R       g709( .A (n298), .B (n339), .C (n964), .Y (n967) );
  NOR2xp33_ASAP7_75t_R      g710( .A (x126), .B (x254), .Y (n968) );
  AND2x2_ASAP7_75t_R        g711( .A (x126), .B (x254), .Y (n969) );
  NOR2xp33_ASAP7_75t_R      g712( .A (n968), .B (n969), .Y (n970) );
  XOR2xp5_ASAP7_75t_R       g713( .A (n967), .B (n970), .Y (y126) );
  MAJIxp5_ASAP7_75t_R       g714( .A (n967), .B (x254), .C (x126), .Y (n972) );
  NOR2xp33_ASAP7_75t_R      g715( .A (x127), .B (x255), .Y (n973) );
  NAND2xp33_ASAP7_75t_R     g716( .A (x127), .B (x255), .Y (n974) );
  INVx1_ASAP7_75t_R         g717( .A (n974), .Y (n975) );
  NOR2xp33_ASAP7_75t_R      g718( .A (n973), .B (n975), .Y (n976) );
  XNOR2xp5_ASAP7_75t_R      g719( .A (n972), .B (n976), .Y (y127) );
  OAI21xp33_ASAP7_75t_R     g720( .A1 (n972), .A2 (n973), .B (n974), .Y (y128) );
endmodule
