module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 ;
  wire n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n281 , n282 , n283 , n284 , n285 , n287 , n288 , n290 , n291 , n292 , n293 , n294 , n296 , n297 , n299 , n300 , n301 , n302 , n303 , n305 , n306 , n308 , n309 , n310 , n311 , n312 , n314 , n315 , n317 , n318 , n319 , n320 , n321 , n323 , n324 , n326 , n327 , n328 , n329 , n330 , n332 , n333 , n334 , n335 , n337 , n338 , n339 , n340 , n341 , n343 , n344 , n345 , n346 , n348 , n349 , n351 , n352 , n354 , n355 , n356 , n357 , n358 , n360 , n361 , n363 , n364 , n366 , n367 , n369 , n370 , n371 , n372 , n373 , n375 , n376 , n378 , n379 , n380 , n381 , n382 , n384 , n385 , n387 , n388 , n389 , n390 , n391 , n393 , n394 , n395 , n396 , n398 , n399 , n401 , n402 , n403 , n404 , n406 , n407 , n408 , n409 , n410 , n412 , n413 , n415 , n416 , n417 , n418 , n419 , n421 , n422 , n423 , n424 , n426 , n427 , n428 , n429 , n430 , n432 , n433 , n434 , n435 , n437 , n438 , n439 , n440 , n441 , n443 , n444 , n445 , n446 , n448 , n449 , n450 , n451 , n452 , n454 , n455 , n457 , n458 , n459 , n460 , n461 , n463 , n464 , n465 , n466 , n468 , n469 , n471 , n472 , n473 , n474 , n476 , n477 , n478 , n479 , n480 , n482 , n483 , n485 , n486 , n487 , n488 , n489 , n491 , n492 , n493 , n494 , n496 , n497 , n499 , n500 , n502 , n503 , n504 , n505 , n506 , n508 , n509 , n511 , n512 , n513 , n514 , n515 , n517 , n518 , n519 , n520 , n522 , n523 , n524 , n525 , n526 , n528 , n529 , n530 , n531 , n533 , n534 , n535 , n536 , n537 , n539 , n540 , n542 , n543 , n545 , n546 , n547 , n548 , n550 , n551 , n552 , n553 , n554 , n556 , n557 , n558 , n559 , n561 , n562 , n563 , n564 , n565 , n567 , n568 , n569 , n570 , n572 , n573 , n574 , n575 , n576 , n578 , n579 , n580 , n581 , n583 , n584 , n585 , n586 , n587 , n589 , n590 , n592 , n593 , n594 , n595 , n596 , n598 , n599 , n600 , n601 , n603 , n604 , n605 , n606 , n607 , n609 , n610 , n611 , n612 , n614 , n615 , n616 , n617 , n618 , n620 , n621 , n623 , n624 , n625 , n626 , n627 , n629 , n630 , n631 , n632 , n634 , n635 , n636 , n637 , n638 , n640 , n641 , n642 , n643 , n645 , n646 , n647 , n648 , n649 , n651 , n652 , n654 , n655 , n656 , n657 , n658 , n660 , n661 , n662 , n663 , n665 , n666 , n667 , n668 , n669 , n671 , n672 , n673 , n674 , n676 , n677 , n678 , n679 , n680 , n682 , n683 , n684 , n685 , n687 , n688 , n690 , n691 , n692 , n693 , n695 , n696 , n697 , n698 , n699 , n701 , n702 , n704 , n705 , n706 , n707 , n708 , n710 , n711 , n713 , n714 , n715 , n716 , n717 , n719 , n720 , n722 , n723 , n724 , n725 , n726 , n728 , n729 , n731 , n732 , n733 , n734 , n735 , n737 , n738 , n739 , n740 , n742 , n743 , n744 , n745 , n746 , n748 , n749 , n751 , n752 , n753 , n754 , n755 , n757 , n758 , n760 , n761 , n762 , n763 , n764 , n766 , n767 , n768 , n769 , n771 , n772 , n774 , n775 , n777 , n778 , n779 , n780 , n781 , n783 , n784 , n785 , n786 , n788 , n789 , n791 , n792 , n793 , n794 , n796 , n797 , n798 , n799 , n800 , n802 , n803 , n805 , n806 , n807 , n808 , n809 , n811 , n812 , n813 , n814 , n816 , n817 , n819 , n820 , n822 , n823 , n824 , n825 , n826 , n828 , n829 , n830 , n831 , n833 , n834 , n835 , n836 , n837 , n839 , n840 , n841 , n842 , n844 , n845 , n846 , n847 , n848 , n850 , n851 , n852 , n853 , n855 , n856 , n857 , n858 , n859 , n861 , n862 , n863 , n864 , n866 , n867 , n868 , n869 , n870 , n872 , n873 , n875 , n876 , n878 , n879 , n880 , n881 , n883 , n884 , n885 , n886 , n887 ;
  XOR2xp5_ASAP7_75t_R    g000( .A (x0), .B (x128), .Y (y0) );
  NAND2xp33_ASAP7_75t_R  g001( .A (x0), .B (x128), .Y (n281) );
  NOR2xp33_ASAP7_75t_R   g002( .A (x1), .B (x129), .Y (n282) );
  INVx1_ASAP7_75t_R      g003( .A (n282), .Y (n283) );
  NAND2xp33_ASAP7_75t_R  g004( .A (x1), .B (x129), .Y (n284) );
  NAND2xp33_ASAP7_75t_R  g005( .A (n283), .B (n284), .Y (n285) );
  XOR2xp5_ASAP7_75t_R    g006( .A (n281), .B (n285), .Y (y1) );
  OAI21xp33_ASAP7_75t_R  g007( .A1 (n282), .A2 (n281), .B (n284), .Y (n287) );
  XOR2xp5_ASAP7_75t_R    g008( .A (x2), .B (x130), .Y (n288) );
  XOR2xp5_ASAP7_75t_R    g009( .A (n287), .B (n288), .Y (y2) );
  MAJIxp5_ASAP7_75t_R    g010( .A (n287), .B (x130), .C (x2), .Y (n290) );
  NOR2xp33_ASAP7_75t_R   g011( .A (x3), .B (x131), .Y (n291) );
  NAND2xp33_ASAP7_75t_R  g012( .A (x3), .B (x131), .Y (n292) );
  INVx1_ASAP7_75t_R      g013( .A (n292), .Y (n293) );
  NOR2xp33_ASAP7_75t_R   g014( .A (n291), .B (n293), .Y (n294) );
  XNOR2xp5_ASAP7_75t_R   g015( .A (n290), .B (n294), .Y (y3) );
  OAI21xp33_ASAP7_75t_R  g016( .A1 (n290), .A2 (n291), .B (n292), .Y (n296) );
  XOR2xp5_ASAP7_75t_R    g017( .A (x4), .B (x132), .Y (n297) );
  XOR2xp5_ASAP7_75t_R    g018( .A (n296), .B (n297), .Y (y4) );
  MAJIxp5_ASAP7_75t_R    g019( .A (n296), .B (x132), .C (x4), .Y (n299) );
  NOR2xp33_ASAP7_75t_R   g020( .A (x5), .B (x133), .Y (n300) );
  NAND2xp33_ASAP7_75t_R  g021( .A (x5), .B (x133), .Y (n301) );
  INVx1_ASAP7_75t_R      g022( .A (n301), .Y (n302) );
  NOR2xp33_ASAP7_75t_R   g023( .A (n300), .B (n302), .Y (n303) );
  XNOR2xp5_ASAP7_75t_R   g024( .A (n299), .B (n303), .Y (y5) );
  OAI21xp33_ASAP7_75t_R  g025( .A1 (n299), .A2 (n300), .B (n301), .Y (n305) );
  XOR2xp5_ASAP7_75t_R    g026( .A (x6), .B (x134), .Y (n306) );
  XOR2xp5_ASAP7_75t_R    g027( .A (n305), .B (n306), .Y (y6) );
  MAJIxp5_ASAP7_75t_R    g028( .A (n305), .B (x134), .C (x6), .Y (n308) );
  NOR2xp33_ASAP7_75t_R   g029( .A (x7), .B (x135), .Y (n309) );
  NAND2xp33_ASAP7_75t_R  g030( .A (x7), .B (x135), .Y (n310) );
  INVx1_ASAP7_75t_R      g031( .A (n310), .Y (n311) );
  NOR2xp33_ASAP7_75t_R   g032( .A (n309), .B (n311), .Y (n312) );
  XNOR2xp5_ASAP7_75t_R   g033( .A (n308), .B (n312), .Y (y7) );
  OAI21xp33_ASAP7_75t_R  g034( .A1 (n308), .A2 (n309), .B (n310), .Y (n314) );
  XOR2xp5_ASAP7_75t_R    g035( .A (x8), .B (x136), .Y (n315) );
  XOR2xp5_ASAP7_75t_R    g036( .A (n314), .B (n315), .Y (y8) );
  MAJIxp5_ASAP7_75t_R    g037( .A (n314), .B (x136), .C (x8), .Y (n317) );
  NOR2xp33_ASAP7_75t_R   g038( .A (x9), .B (x137), .Y (n318) );
  NAND2xp33_ASAP7_75t_R  g039( .A (x9), .B (x137), .Y (n319) );
  INVx1_ASAP7_75t_R      g040( .A (n319), .Y (n320) );
  NOR2xp33_ASAP7_75t_R   g041( .A (n318), .B (n320), .Y (n321) );
  XNOR2xp5_ASAP7_75t_R   g042( .A (n317), .B (n321), .Y (y9) );
  OAI21xp33_ASAP7_75t_R  g043( .A1 (n317), .A2 (n318), .B (n319), .Y (n323) );
  XOR2xp5_ASAP7_75t_R    g044( .A (x10), .B (x138), .Y (n324) );
  XOR2xp5_ASAP7_75t_R    g045( .A (n323), .B (n324), .Y (y10) );
  NOR2xp33_ASAP7_75t_R   g046( .A (x11), .B (x139), .Y (n327) );
  INVx1_ASAP7_75t_R      g047( .A (n327), .Y (n328) );
  NAND2xp33_ASAP7_75t_R  g048( .A (x11), .B (x139), .Y (n329) );
  NAND2xp33_ASAP7_75t_R  g049( .A (n328), .B (n329), .Y (n330) );
  MAJIxp5_ASAP7_75t_R    g050( .A (n323), .B (x138), .C (x10), .Y (n326) );
  XOR2xp5_ASAP7_75t_R    g051( .A (n330), .B (n326), .Y (y11) );
  OAI21xp33_ASAP7_75t_R  g052( .A1 (n326), .A2 (n327), .B (n329), .Y (n332) );
  NOR2xp33_ASAP7_75t_R   g053( .A (x12), .B (x140), .Y (n333) );
  AND2x2_ASAP7_75t_R     g054( .A (x12), .B (x140), .Y (n334) );
  NOR2xp33_ASAP7_75t_R   g055( .A (n333), .B (n334), .Y (n335) );
  XOR2xp5_ASAP7_75t_R    g056( .A (n332), .B (n335), .Y (y12) );
  MAJIxp5_ASAP7_75t_R    g057( .A (n332), .B (x140), .C (x12), .Y (n337) );
  NOR2xp33_ASAP7_75t_R   g058( .A (x13), .B (x141), .Y (n338) );
  NAND2xp33_ASAP7_75t_R  g059( .A (x13), .B (x141), .Y (n339) );
  INVx1_ASAP7_75t_R      g060( .A (n339), .Y (n340) );
  NOR2xp33_ASAP7_75t_R   g061( .A (n338), .B (n340), .Y (n341) );
  XNOR2xp5_ASAP7_75t_R   g062( .A (n337), .B (n341), .Y (y13) );
  OAI21xp33_ASAP7_75t_R  g063( .A1 (n337), .A2 (n338), .B (n339), .Y (n343) );
  NOR2xp33_ASAP7_75t_R   g064( .A (x14), .B (x142), .Y (n344) );
  AND2x2_ASAP7_75t_R     g065( .A (x14), .B (x142), .Y (n345) );
  NOR2xp33_ASAP7_75t_R   g066( .A (n344), .B (n345), .Y (n346) );
  XOR2xp5_ASAP7_75t_R    g067( .A (n343), .B (n346), .Y (y14) );
  MAJIxp5_ASAP7_75t_R    g068( .A (n343), .B (x142), .C (x14), .Y (n348) );
  XOR2xp5_ASAP7_75t_R    g069( .A (x15), .B (x143), .Y (n349) );
  XNOR2xp5_ASAP7_75t_R   g070( .A (n348), .B (n349), .Y (y15) );
  INVx1_ASAP7_75t_R      g071( .A (x15), .Y (n258) );
  INVx1_ASAP7_75t_R      g072( .A (x143), .Y (n269) );
  MAJIxp5_ASAP7_75t_R    g073( .A (n258), .B (n269), .C (n348), .Y (n351) );
  XOR2xp5_ASAP7_75t_R    g074( .A (x16), .B (x144), .Y (n352) );
  XOR2xp5_ASAP7_75t_R    g075( .A (n351), .B (n352), .Y (y16) );
  NOR2xp33_ASAP7_75t_R   g076( .A (x17), .B (x145), .Y (n355) );
  INVx1_ASAP7_75t_R      g077( .A (n355), .Y (n356) );
  NAND2xp33_ASAP7_75t_R  g078( .A (x17), .B (x145), .Y (n357) );
  NAND2xp33_ASAP7_75t_R  g079( .A (n356), .B (n357), .Y (n358) );
  MAJIxp5_ASAP7_75t_R    g080( .A (n351), .B (x144), .C (x16), .Y (n354) );
  XOR2xp5_ASAP7_75t_R    g081( .A (n358), .B (n354), .Y (y17) );
  OAI21xp33_ASAP7_75t_R  g082( .A1 (n354), .A2 (n355), .B (n357), .Y (n360) );
  XOR2xp5_ASAP7_75t_R    g083( .A (x18), .B (x146), .Y (n361) );
  XOR2xp5_ASAP7_75t_R    g084( .A (n360), .B (n361), .Y (y18) );
  MAJIxp5_ASAP7_75t_R    g085( .A (n360), .B (x146), .C (x18), .Y (n363) );
  XOR2xp5_ASAP7_75t_R    g086( .A (x19), .B (x147), .Y (n364) );
  XNOR2xp5_ASAP7_75t_R   g087( .A (n363), .B (n364), .Y (y19) );
  INVx1_ASAP7_75t_R      g088( .A (x19), .Y (n259) );
  INVx1_ASAP7_75t_R      g089( .A (x147), .Y (n270) );
  MAJIxp5_ASAP7_75t_R    g090( .A (n259), .B (n270), .C (n363), .Y (n366) );
  XOR2xp5_ASAP7_75t_R    g091( .A (x20), .B (x148), .Y (n367) );
  XOR2xp5_ASAP7_75t_R    g092( .A (n366), .B (n367), .Y (y20) );
  NOR2xp33_ASAP7_75t_R   g093( .A (x21), .B (x149), .Y (n370) );
  INVx1_ASAP7_75t_R      g094( .A (n370), .Y (n371) );
  NAND2xp33_ASAP7_75t_R  g095( .A (x21), .B (x149), .Y (n372) );
  NAND2xp33_ASAP7_75t_R  g096( .A (n371), .B (n372), .Y (n373) );
  MAJIxp5_ASAP7_75t_R    g097( .A (n366), .B (x148), .C (x20), .Y (n369) );
  XOR2xp5_ASAP7_75t_R    g098( .A (n373), .B (n369), .Y (y21) );
  OAI21xp33_ASAP7_75t_R  g099( .A1 (n369), .A2 (n370), .B (n372), .Y (n375) );
  XOR2xp5_ASAP7_75t_R    g100( .A (x22), .B (x150), .Y (n376) );
  XOR2xp5_ASAP7_75t_R    g101( .A (n375), .B (n376), .Y (y22) );
  MAJIxp5_ASAP7_75t_R    g102( .A (n375), .B (x150), .C (x22), .Y (n378) );
  NOR2xp33_ASAP7_75t_R   g103( .A (x23), .B (x151), .Y (n379) );
  NAND2xp33_ASAP7_75t_R  g104( .A (x23), .B (x151), .Y (n380) );
  INVx1_ASAP7_75t_R      g105( .A (n380), .Y (n381) );
  NOR2xp33_ASAP7_75t_R   g106( .A (n379), .B (n381), .Y (n382) );
  XNOR2xp5_ASAP7_75t_R   g107( .A (n378), .B (n382), .Y (y23) );
  OAI21xp33_ASAP7_75t_R  g108( .A1 (n378), .A2 (n379), .B (n380), .Y (n384) );
  XNOR2xp5_ASAP7_75t_R   g109( .A (x24), .B (x152), .Y (n385) );
  XNOR2xp5_ASAP7_75t_R   g110( .A (n384), .B (n385), .Y (y24) );
  MAJIxp5_ASAP7_75t_R    g111( .A (n384), .B (x152), .C (x24), .Y (n387) );
  NOR2xp33_ASAP7_75t_R   g112( .A (x25), .B (x153), .Y (n388) );
  NAND2xp33_ASAP7_75t_R  g113( .A (x25), .B (x153), .Y (n389) );
  INVx1_ASAP7_75t_R      g114( .A (n389), .Y (n390) );
  NOR2xp33_ASAP7_75t_R   g115( .A (n388), .B (n390), .Y (n391) );
  XNOR2xp5_ASAP7_75t_R   g116( .A (n387), .B (n391), .Y (y25) );
  OAI21xp33_ASAP7_75t_R  g117( .A1 (n387), .A2 (n388), .B (n389), .Y (n393) );
  NOR2xp33_ASAP7_75t_R   g118( .A (x26), .B (x154), .Y (n394) );
  AND2x2_ASAP7_75t_R     g119( .A (x26), .B (x154), .Y (n395) );
  NOR2xp33_ASAP7_75t_R   g120( .A (n394), .B (n395), .Y (n396) );
  XOR2xp5_ASAP7_75t_R    g121( .A (n393), .B (n396), .Y (y26) );
  MAJIxp5_ASAP7_75t_R    g122( .A (n393), .B (x154), .C (x26), .Y (n398) );
  XOR2xp5_ASAP7_75t_R    g123( .A (x27), .B (x155), .Y (n399) );
  XNOR2xp5_ASAP7_75t_R   g124( .A (n398), .B (n399), .Y (y27) );
  INVx1_ASAP7_75t_R      g125( .A (x27), .Y (n260) );
  INVx1_ASAP7_75t_R      g126( .A (x155), .Y (n271) );
  MAJIxp5_ASAP7_75t_R    g127( .A (n260), .B (n271), .C (n398), .Y (n401) );
  OR2x2_ASAP7_75t_R      g128( .A (x28), .B (x156), .Y (n402) );
  NAND2xp33_ASAP7_75t_R  g129( .A (x28), .B (x156), .Y (n403) );
  NAND2xp33_ASAP7_75t_R  g130( .A (n402), .B (n403), .Y (n404) );
  XNOR2xp5_ASAP7_75t_R   g131( .A (n401), .B (n404), .Y (y28) );
  NOR2xp33_ASAP7_75t_R   g132( .A (x29), .B (x157), .Y (n407) );
  INVx1_ASAP7_75t_R      g133( .A (n407), .Y (n408) );
  NAND2xp33_ASAP7_75t_R  g134( .A (x29), .B (x157), .Y (n409) );
  NAND2xp33_ASAP7_75t_R  g135( .A (n408), .B (n409), .Y (n410) );
  MAJIxp5_ASAP7_75t_R    g136( .A (n401), .B (x156), .C (x28), .Y (n406) );
  XOR2xp5_ASAP7_75t_R    g137( .A (n410), .B (n406), .Y (y29) );
  OAI21xp33_ASAP7_75t_R  g138( .A1 (n406), .A2 (n407), .B (n409), .Y (n412) );
  XOR2xp5_ASAP7_75t_R    g139( .A (x30), .B (x158), .Y (n413) );
  XOR2xp5_ASAP7_75t_R    g140( .A (n412), .B (n413), .Y (y30) );
  NOR2xp33_ASAP7_75t_R   g141( .A (x31), .B (x159), .Y (n416) );
  INVx1_ASAP7_75t_R      g142( .A (n416), .Y (n417) );
  NAND2xp33_ASAP7_75t_R  g143( .A (x31), .B (x159), .Y (n418) );
  NAND2xp33_ASAP7_75t_R  g144( .A (n417), .B (n418), .Y (n419) );
  MAJIxp5_ASAP7_75t_R    g145( .A (n412), .B (x158), .C (x30), .Y (n415) );
  XOR2xp5_ASAP7_75t_R    g146( .A (n419), .B (n415), .Y (y31) );
  OAI21xp33_ASAP7_75t_R  g147( .A1 (n415), .A2 (n416), .B (n418), .Y (n421) );
  NOR2xp33_ASAP7_75t_R   g148( .A (x32), .B (x160), .Y (n422) );
  AND2x2_ASAP7_75t_R     g149( .A (x32), .B (x160), .Y (n423) );
  NOR2xp33_ASAP7_75t_R   g150( .A (n422), .B (n423), .Y (n424) );
  XOR2xp5_ASAP7_75t_R    g151( .A (n421), .B (n424), .Y (y32) );
  MAJIxp5_ASAP7_75t_R    g152( .A (n421), .B (x160), .C (x32), .Y (n426) );
  NOR2xp33_ASAP7_75t_R   g153( .A (x33), .B (x161), .Y (n427) );
  NAND2xp33_ASAP7_75t_R  g154( .A (x33), .B (x161), .Y (n428) );
  INVx1_ASAP7_75t_R      g155( .A (n428), .Y (n429) );
  NOR2xp33_ASAP7_75t_R   g156( .A (n427), .B (n429), .Y (n430) );
  XNOR2xp5_ASAP7_75t_R   g157( .A (n426), .B (n430), .Y (y33) );
  OAI21xp33_ASAP7_75t_R  g158( .A1 (n426), .A2 (n427), .B (n428), .Y (n432) );
  OR2x2_ASAP7_75t_R      g159( .A (x34), .B (x162), .Y (n433) );
  NAND2xp33_ASAP7_75t_R  g160( .A (x34), .B (x162), .Y (n434) );
  NAND2xp33_ASAP7_75t_R  g161( .A (n433), .B (n434), .Y (n435) );
  XNOR2xp5_ASAP7_75t_R   g162( .A (n432), .B (n435), .Y (y34) );
  NOR2xp33_ASAP7_75t_R   g163( .A (x35), .B (x163), .Y (n438) );
  INVx1_ASAP7_75t_R      g164( .A (n438), .Y (n439) );
  NAND2xp33_ASAP7_75t_R  g165( .A (x35), .B (x163), .Y (n440) );
  NAND2xp33_ASAP7_75t_R  g166( .A (n439), .B (n440), .Y (n441) );
  MAJIxp5_ASAP7_75t_R    g167( .A (n432), .B (x162), .C (x34), .Y (n437) );
  XOR2xp5_ASAP7_75t_R    g168( .A (n441), .B (n437), .Y (y35) );
  OAI21xp33_ASAP7_75t_R  g169( .A1 (n437), .A2 (n438), .B (n440), .Y (n443) );
  NOR2xp33_ASAP7_75t_R   g170( .A (x36), .B (x164), .Y (n444) );
  AND2x2_ASAP7_75t_R     g171( .A (x36), .B (x164), .Y (n445) );
  NOR2xp33_ASAP7_75t_R   g172( .A (n444), .B (n445), .Y (n446) );
  XOR2xp5_ASAP7_75t_R    g173( .A (n443), .B (n446), .Y (y36) );
  MAJIxp5_ASAP7_75t_R    g174( .A (n443), .B (x164), .C (x36), .Y (n448) );
  NOR2xp33_ASAP7_75t_R   g175( .A (x37), .B (x165), .Y (n449) );
  NAND2xp33_ASAP7_75t_R  g176( .A (x37), .B (x165), .Y (n450) );
  INVx1_ASAP7_75t_R      g177( .A (n450), .Y (n451) );
  NOR2xp33_ASAP7_75t_R   g178( .A (n449), .B (n451), .Y (n452) );
  XNOR2xp5_ASAP7_75t_R   g179( .A (n448), .B (n452), .Y (y37) );
  OAI21xp33_ASAP7_75t_R  g180( .A1 (n448), .A2 (n449), .B (n450), .Y (n454) );
  XNOR2xp5_ASAP7_75t_R   g181( .A (x38), .B (x166), .Y (n455) );
  XNOR2xp5_ASAP7_75t_R   g182( .A (n454), .B (n455), .Y (y38) );
  NOR2xp33_ASAP7_75t_R   g183( .A (x39), .B (x167), .Y (n458) );
  INVx1_ASAP7_75t_R      g184( .A (n458), .Y (n459) );
  NAND2xp33_ASAP7_75t_R  g185( .A (x39), .B (x167), .Y (n460) );
  NAND2xp33_ASAP7_75t_R  g186( .A (n459), .B (n460), .Y (n461) );
  MAJIxp5_ASAP7_75t_R    g187( .A (n454), .B (x166), .C (x38), .Y (n457) );
  XOR2xp5_ASAP7_75t_R    g188( .A (n461), .B (n457), .Y (y39) );
  OAI21xp33_ASAP7_75t_R  g189( .A1 (n457), .A2 (n458), .B (n460), .Y (n463) );
  NOR2xp33_ASAP7_75t_R   g190( .A (x40), .B (x168), .Y (n464) );
  AND2x2_ASAP7_75t_R     g191( .A (x40), .B (x168), .Y (n465) );
  NOR2xp33_ASAP7_75t_R   g192( .A (n464), .B (n465), .Y (n466) );
  XOR2xp5_ASAP7_75t_R    g193( .A (n463), .B (n466), .Y (y40) );
  MAJIxp5_ASAP7_75t_R    g194( .A (n463), .B (x168), .C (x40), .Y (n468) );
  XOR2xp5_ASAP7_75t_R    g195( .A (x41), .B (x169), .Y (n469) );
  XNOR2xp5_ASAP7_75t_R   g196( .A (n468), .B (n469), .Y (y41) );
  INVx1_ASAP7_75t_R      g197( .A (x41), .Y (n261) );
  INVx1_ASAP7_75t_R      g198( .A (x169), .Y (n272) );
  MAJIxp5_ASAP7_75t_R    g199( .A (n261), .B (n272), .C (n468), .Y (n471) );
  OR2x2_ASAP7_75t_R      g200( .A (x42), .B (x170), .Y (n472) );
  NAND2xp33_ASAP7_75t_R  g201( .A (x42), .B (x170), .Y (n473) );
  NAND2xp33_ASAP7_75t_R  g202( .A (n472), .B (n473), .Y (n474) );
  XNOR2xp5_ASAP7_75t_R   g203( .A (n471), .B (n474), .Y (y42) );
  NOR2xp33_ASAP7_75t_R   g204( .A (x43), .B (x171), .Y (n477) );
  INVx1_ASAP7_75t_R      g205( .A (n477), .Y (n478) );
  NAND2xp33_ASAP7_75t_R  g206( .A (x43), .B (x171), .Y (n479) );
  NAND2xp33_ASAP7_75t_R  g207( .A (n478), .B (n479), .Y (n480) );
  MAJIxp5_ASAP7_75t_R    g208( .A (n471), .B (x170), .C (x42), .Y (n476) );
  XOR2xp5_ASAP7_75t_R    g209( .A (n480), .B (n476), .Y (y43) );
  OAI21xp33_ASAP7_75t_R  g210( .A1 (n476), .A2 (n477), .B (n479), .Y (n482) );
  XOR2xp5_ASAP7_75t_R    g211( .A (x44), .B (x172), .Y (n483) );
  XOR2xp5_ASAP7_75t_R    g212( .A (n482), .B (n483), .Y (y44) );
  MAJIxp5_ASAP7_75t_R    g213( .A (n482), .B (x172), .C (x44), .Y (n485) );
  NOR2xp33_ASAP7_75t_R   g214( .A (x45), .B (x173), .Y (n486) );
  NAND2xp33_ASAP7_75t_R  g215( .A (x45), .B (x173), .Y (n487) );
  INVx1_ASAP7_75t_R      g216( .A (n487), .Y (n488) );
  NOR2xp33_ASAP7_75t_R   g217( .A (n486), .B (n488), .Y (n489) );
  XNOR2xp5_ASAP7_75t_R   g218( .A (n485), .B (n489), .Y (y45) );
  OAI21xp33_ASAP7_75t_R  g219( .A1 (n485), .A2 (n486), .B (n487), .Y (n491) );
  NOR2xp33_ASAP7_75t_R   g220( .A (x46), .B (x174), .Y (n492) );
  AND2x2_ASAP7_75t_R     g221( .A (x46), .B (x174), .Y (n493) );
  NOR2xp33_ASAP7_75t_R   g222( .A (n492), .B (n493), .Y (n494) );
  XOR2xp5_ASAP7_75t_R    g223( .A (n491), .B (n494), .Y (y46) );
  MAJIxp5_ASAP7_75t_R    g224( .A (n491), .B (x174), .C (x46), .Y (n496) );
  XOR2xp5_ASAP7_75t_R    g225( .A (x47), .B (x175), .Y (n497) );
  XNOR2xp5_ASAP7_75t_R   g226( .A (n496), .B (n497), .Y (y47) );
  INVx1_ASAP7_75t_R      g227( .A (x47), .Y (n262) );
  INVx1_ASAP7_75t_R      g228( .A (x175), .Y (n273) );
  MAJIxp5_ASAP7_75t_R    g229( .A (n262), .B (n273), .C (n496), .Y (n499) );
  XOR2xp5_ASAP7_75t_R    g230( .A (x48), .B (x176), .Y (n500) );
  XOR2xp5_ASAP7_75t_R    g231( .A (n499), .B (n500), .Y (y48) );
  NOR2xp33_ASAP7_75t_R   g232( .A (x49), .B (x177), .Y (n503) );
  INVx1_ASAP7_75t_R      g233( .A (n503), .Y (n504) );
  NAND2xp33_ASAP7_75t_R  g234( .A (x49), .B (x177), .Y (n505) );
  NAND2xp33_ASAP7_75t_R  g235( .A (n504), .B (n505), .Y (n506) );
  MAJIxp5_ASAP7_75t_R    g236( .A (n499), .B (x176), .C (x48), .Y (n502) );
  XOR2xp5_ASAP7_75t_R    g237( .A (n506), .B (n502), .Y (y49) );
  OAI21xp33_ASAP7_75t_R  g238( .A1 (n502), .A2 (n503), .B (n505), .Y (n508) );
  XOR2xp5_ASAP7_75t_R    g239( .A (x50), .B (x178), .Y (n509) );
  XOR2xp5_ASAP7_75t_R    g240( .A (n508), .B (n509), .Y (y50) );
  MAJIxp5_ASAP7_75t_R    g241( .A (n508), .B (x178), .C (x50), .Y (n511) );
  NOR2xp33_ASAP7_75t_R   g242( .A (x51), .B (x179), .Y (n512) );
  NAND2xp33_ASAP7_75t_R  g243( .A (x51), .B (x179), .Y (n513) );
  INVx1_ASAP7_75t_R      g244( .A (n513), .Y (n514) );
  NOR2xp33_ASAP7_75t_R   g245( .A (n512), .B (n514), .Y (n515) );
  XNOR2xp5_ASAP7_75t_R   g246( .A (n511), .B (n515), .Y (y51) );
  OAI21xp33_ASAP7_75t_R  g247( .A1 (n511), .A2 (n512), .B (n513), .Y (n517) );
  NOR2xp33_ASAP7_75t_R   g248( .A (x52), .B (x180), .Y (n518) );
  AND2x2_ASAP7_75t_R     g249( .A (x52), .B (x180), .Y (n519) );
  NOR2xp33_ASAP7_75t_R   g250( .A (n518), .B (n519), .Y (n520) );
  XOR2xp5_ASAP7_75t_R    g251( .A (n517), .B (n520), .Y (y52) );
  MAJIxp5_ASAP7_75t_R    g252( .A (n517), .B (x180), .C (x52), .Y (n522) );
  NOR2xp33_ASAP7_75t_R   g253( .A (x53), .B (x181), .Y (n523) );
  NAND2xp33_ASAP7_75t_R  g254( .A (x53), .B (x181), .Y (n524) );
  INVx1_ASAP7_75t_R      g255( .A (n524), .Y (n525) );
  NOR2xp33_ASAP7_75t_R   g256( .A (n523), .B (n525), .Y (n526) );
  XNOR2xp5_ASAP7_75t_R   g257( .A (n522), .B (n526), .Y (y53) );
  OAI21xp33_ASAP7_75t_R  g258( .A1 (n522), .A2 (n523), .B (n524), .Y (n528) );
  NOR2xp33_ASAP7_75t_R   g259( .A (x54), .B (x182), .Y (n529) );
  AND2x2_ASAP7_75t_R     g260( .A (x54), .B (x182), .Y (n530) );
  NOR2xp33_ASAP7_75t_R   g261( .A (n529), .B (n530), .Y (n531) );
  XOR2xp5_ASAP7_75t_R    g262( .A (n528), .B (n531), .Y (y54) );
  MAJIxp5_ASAP7_75t_R    g263( .A (n528), .B (x182), .C (x54), .Y (n533) );
  NOR2xp33_ASAP7_75t_R   g264( .A (x55), .B (x183), .Y (n534) );
  NAND2xp33_ASAP7_75t_R  g265( .A (x55), .B (x183), .Y (n535) );
  INVx1_ASAP7_75t_R      g266( .A (n535), .Y (n536) );
  NOR2xp33_ASAP7_75t_R   g267( .A (n534), .B (n536), .Y (n537) );
  XNOR2xp5_ASAP7_75t_R   g268( .A (n533), .B (n537), .Y (y55) );
  OAI21xp33_ASAP7_75t_R  g269( .A1 (n533), .A2 (n534), .B (n535), .Y (n539) );
  XOR2xp5_ASAP7_75t_R    g270( .A (x56), .B (x184), .Y (n540) );
  XOR2xp5_ASAP7_75t_R    g271( .A (n539), .B (n540), .Y (y56) );
  MAJIxp5_ASAP7_75t_R    g272( .A (n539), .B (x184), .C (x56), .Y (n542) );
  XOR2xp5_ASAP7_75t_R    g273( .A (x57), .B (x185), .Y (n543) );
  XNOR2xp5_ASAP7_75t_R   g274( .A (n542), .B (n543), .Y (y57) );
  INVx1_ASAP7_75t_R      g275( .A (x57), .Y (n263) );
  INVx1_ASAP7_75t_R      g276( .A (x185), .Y (n274) );
  MAJIxp5_ASAP7_75t_R    g277( .A (n263), .B (n274), .C (n542), .Y (n545) );
  OR2x2_ASAP7_75t_R      g278( .A (x58), .B (x186), .Y (n546) );
  NAND2xp33_ASAP7_75t_R  g279( .A (x58), .B (x186), .Y (n547) );
  NAND2xp33_ASAP7_75t_R  g280( .A (n546), .B (n547), .Y (n548) );
  XNOR2xp5_ASAP7_75t_R   g281( .A (n545), .B (n548), .Y (y58) );
  NOR2xp33_ASAP7_75t_R   g282( .A (x59), .B (x187), .Y (n551) );
  INVx1_ASAP7_75t_R      g283( .A (n551), .Y (n552) );
  NAND2xp33_ASAP7_75t_R  g284( .A (x59), .B (x187), .Y (n553) );
  NAND2xp33_ASAP7_75t_R  g285( .A (n552), .B (n553), .Y (n554) );
  MAJIxp5_ASAP7_75t_R    g286( .A (n545), .B (x186), .C (x58), .Y (n550) );
  XOR2xp5_ASAP7_75t_R    g287( .A (n554), .B (n550), .Y (y59) );
  OAI21xp33_ASAP7_75t_R  g288( .A1 (n550), .A2 (n551), .B (n553), .Y (n556) );
  NOR2xp33_ASAP7_75t_R   g289( .A (x60), .B (x188), .Y (n557) );
  AND2x2_ASAP7_75t_R     g290( .A (x60), .B (x188), .Y (n558) );
  NOR2xp33_ASAP7_75t_R   g291( .A (n557), .B (n558), .Y (n559) );
  XOR2xp5_ASAP7_75t_R    g292( .A (n556), .B (n559), .Y (y60) );
  MAJIxp5_ASAP7_75t_R    g293( .A (n556), .B (x188), .C (x60), .Y (n561) );
  NOR2xp33_ASAP7_75t_R   g294( .A (x61), .B (x189), .Y (n562) );
  NAND2xp33_ASAP7_75t_R  g295( .A (x61), .B (x189), .Y (n563) );
  INVx1_ASAP7_75t_R      g296( .A (n563), .Y (n564) );
  NOR2xp33_ASAP7_75t_R   g297( .A (n562), .B (n564), .Y (n565) );
  XNOR2xp5_ASAP7_75t_R   g298( .A (n561), .B (n565), .Y (y61) );
  OAI21xp33_ASAP7_75t_R  g299( .A1 (n561), .A2 (n562), .B (n563), .Y (n567) );
  NOR2xp33_ASAP7_75t_R   g300( .A (x62), .B (x190), .Y (n568) );
  AND2x2_ASAP7_75t_R     g301( .A (x62), .B (x190), .Y (n569) );
  NOR2xp33_ASAP7_75t_R   g302( .A (n568), .B (n569), .Y (n570) );
  XOR2xp5_ASAP7_75t_R    g303( .A (n567), .B (n570), .Y (y62) );
  MAJIxp5_ASAP7_75t_R    g304( .A (n567), .B (x190), .C (x62), .Y (n572) );
  NOR2xp33_ASAP7_75t_R   g305( .A (x63), .B (x191), .Y (n573) );
  NAND2xp33_ASAP7_75t_R  g306( .A (x63), .B (x191), .Y (n574) );
  INVx1_ASAP7_75t_R      g307( .A (n574), .Y (n575) );
  NOR2xp33_ASAP7_75t_R   g308( .A (n573), .B (n575), .Y (n576) );
  XNOR2xp5_ASAP7_75t_R   g309( .A (n572), .B (n576), .Y (y63) );
  OAI21xp33_ASAP7_75t_R  g310( .A1 (n572), .A2 (n573), .B (n574), .Y (n578) );
  NOR2xp33_ASAP7_75t_R   g311( .A (x64), .B (x192), .Y (n579) );
  AND2x2_ASAP7_75t_R     g312( .A (x64), .B (x192), .Y (n580) );
  NOR2xp33_ASAP7_75t_R   g313( .A (n579), .B (n580), .Y (n581) );
  XOR2xp5_ASAP7_75t_R    g314( .A (n578), .B (n581), .Y (y64) );
  MAJIxp5_ASAP7_75t_R    g315( .A (n578), .B (x192), .C (x64), .Y (n583) );
  NOR2xp33_ASAP7_75t_R   g316( .A (x65), .B (x193), .Y (n584) );
  NAND2xp33_ASAP7_75t_R  g317( .A (x65), .B (x193), .Y (n585) );
  INVx1_ASAP7_75t_R      g318( .A (n585), .Y (n586) );
  NOR2xp33_ASAP7_75t_R   g319( .A (n584), .B (n586), .Y (n587) );
  XNOR2xp5_ASAP7_75t_R   g320( .A (n583), .B (n587), .Y (y65) );
  OAI21xp33_ASAP7_75t_R  g321( .A1 (n583), .A2 (n584), .B (n585), .Y (n589) );
  XOR2xp5_ASAP7_75t_R    g322( .A (x66), .B (x194), .Y (n590) );
  XOR2xp5_ASAP7_75t_R    g323( .A (n589), .B (n590), .Y (y66) );
  MAJIxp5_ASAP7_75t_R    g324( .A (n589), .B (x194), .C (x66), .Y (n592) );
  NOR2xp33_ASAP7_75t_R   g325( .A (x67), .B (x195), .Y (n593) );
  NAND2xp33_ASAP7_75t_R  g326( .A (x67), .B (x195), .Y (n594) );
  INVx1_ASAP7_75t_R      g327( .A (n594), .Y (n595) );
  NOR2xp33_ASAP7_75t_R   g328( .A (n593), .B (n595), .Y (n596) );
  XNOR2xp5_ASAP7_75t_R   g329( .A (n592), .B (n596), .Y (y67) );
  OAI21xp33_ASAP7_75t_R  g330( .A1 (n592), .A2 (n593), .B (n594), .Y (n598) );
  NOR2xp33_ASAP7_75t_R   g331( .A (x68), .B (x196), .Y (n599) );
  AND2x2_ASAP7_75t_R     g332( .A (x68), .B (x196), .Y (n600) );
  NOR2xp33_ASAP7_75t_R   g333( .A (n599), .B (n600), .Y (n601) );
  XOR2xp5_ASAP7_75t_R    g334( .A (n598), .B (n601), .Y (y68) );
  MAJIxp5_ASAP7_75t_R    g335( .A (n598), .B (x196), .C (x68), .Y (n603) );
  NOR2xp33_ASAP7_75t_R   g336( .A (x69), .B (x197), .Y (n604) );
  NAND2xp33_ASAP7_75t_R  g337( .A (x69), .B (x197), .Y (n605) );
  INVx1_ASAP7_75t_R      g338( .A (n605), .Y (n606) );
  NOR2xp33_ASAP7_75t_R   g339( .A (n604), .B (n606), .Y (n607) );
  XNOR2xp5_ASAP7_75t_R   g340( .A (n603), .B (n607), .Y (y69) );
  OAI21xp33_ASAP7_75t_R  g341( .A1 (n603), .A2 (n604), .B (n605), .Y (n609) );
  OR2x2_ASAP7_75t_R      g342( .A (x70), .B (x198), .Y (n610) );
  NAND2xp33_ASAP7_75t_R  g343( .A (x70), .B (x198), .Y (n611) );
  NAND2xp33_ASAP7_75t_R  g344( .A (n610), .B (n611), .Y (n612) );
  XNOR2xp5_ASAP7_75t_R   g345( .A (n609), .B (n612), .Y (y70) );
  MAJIxp5_ASAP7_75t_R    g346( .A (n609), .B (x198), .C (x70), .Y (n614) );
  NOR2xp33_ASAP7_75t_R   g347( .A (x71), .B (x199), .Y (n615) );
  NAND2xp33_ASAP7_75t_R  g348( .A (x71), .B (x199), .Y (n616) );
  INVx1_ASAP7_75t_R      g349( .A (n616), .Y (n617) );
  NOR2xp33_ASAP7_75t_R   g350( .A (n615), .B (n617), .Y (n618) );
  XNOR2xp5_ASAP7_75t_R   g351( .A (n614), .B (n618), .Y (y71) );
  OAI21xp33_ASAP7_75t_R  g352( .A1 (n614), .A2 (n615), .B (n616), .Y (n620) );
  XOR2xp5_ASAP7_75t_R    g353( .A (x72), .B (x200), .Y (n621) );
  XOR2xp5_ASAP7_75t_R    g354( .A (n620), .B (n621), .Y (y72) );
  MAJIxp5_ASAP7_75t_R    g355( .A (n620), .B (x200), .C (x72), .Y (n623) );
  NOR2xp33_ASAP7_75t_R   g356( .A (x73), .B (x201), .Y (n624) );
  NAND2xp33_ASAP7_75t_R  g357( .A (x73), .B (x201), .Y (n625) );
  INVx1_ASAP7_75t_R      g358( .A (n625), .Y (n626) );
  NOR2xp33_ASAP7_75t_R   g359( .A (n624), .B (n626), .Y (n627) );
  XNOR2xp5_ASAP7_75t_R   g360( .A (n623), .B (n627), .Y (y73) );
  OAI21xp33_ASAP7_75t_R  g361( .A1 (n623), .A2 (n624), .B (n625), .Y (n629) );
  NOR2xp33_ASAP7_75t_R   g362( .A (x74), .B (x202), .Y (n630) );
  AND2x2_ASAP7_75t_R     g363( .A (x74), .B (x202), .Y (n631) );
  NOR2xp33_ASAP7_75t_R   g364( .A (n630), .B (n631), .Y (n632) );
  XOR2xp5_ASAP7_75t_R    g365( .A (n629), .B (n632), .Y (y74) );
  MAJIxp5_ASAP7_75t_R    g366( .A (n629), .B (x202), .C (x74), .Y (n634) );
  NOR2xp33_ASAP7_75t_R   g367( .A (x75), .B (x203), .Y (n635) );
  NAND2xp33_ASAP7_75t_R  g368( .A (x75), .B (x203), .Y (n636) );
  INVx1_ASAP7_75t_R      g369( .A (n636), .Y (n637) );
  NOR2xp33_ASAP7_75t_R   g370( .A (n635), .B (n637), .Y (n638) );
  XNOR2xp5_ASAP7_75t_R   g371( .A (n634), .B (n638), .Y (y75) );
  OAI21xp33_ASAP7_75t_R  g372( .A1 (n634), .A2 (n635), .B (n636), .Y (n640) );
  OR2x2_ASAP7_75t_R      g373( .A (x76), .B (x204), .Y (n641) );
  NAND2xp33_ASAP7_75t_R  g374( .A (x76), .B (x204), .Y (n642) );
  AND2x2_ASAP7_75t_R     g375( .A (n641), .B (n642), .Y (n643) );
  XOR2xp5_ASAP7_75t_R    g376( .A (n640), .B (n643), .Y (y76) );
  MAJIxp5_ASAP7_75t_R    g377( .A (n640), .B (x204), .C (x76), .Y (n645) );
  NOR2xp33_ASAP7_75t_R   g378( .A (x77), .B (x205), .Y (n646) );
  NAND2xp33_ASAP7_75t_R  g379( .A (x77), .B (x205), .Y (n647) );
  INVx1_ASAP7_75t_R      g380( .A (n647), .Y (n648) );
  NOR2xp33_ASAP7_75t_R   g381( .A (n646), .B (n648), .Y (n649) );
  XNOR2xp5_ASAP7_75t_R   g382( .A (n645), .B (n649), .Y (y77) );
  OAI21xp33_ASAP7_75t_R  g383( .A1 (n645), .A2 (n646), .B (n647), .Y (n651) );
  XNOR2xp5_ASAP7_75t_R   g384( .A (x78), .B (x206), .Y (n652) );
  XNOR2xp5_ASAP7_75t_R   g385( .A (n651), .B (n652), .Y (y78) );
  NOR2xp33_ASAP7_75t_R   g386( .A (x79), .B (x207), .Y (n655) );
  INVx1_ASAP7_75t_R      g387( .A (n655), .Y (n656) );
  NAND2xp33_ASAP7_75t_R  g388( .A (x79), .B (x207), .Y (n657) );
  NAND2xp33_ASAP7_75t_R  g389( .A (n656), .B (n657), .Y (n658) );
  MAJIxp5_ASAP7_75t_R    g390( .A (n651), .B (x206), .C (x78), .Y (n654) );
  XOR2xp5_ASAP7_75t_R    g391( .A (n658), .B (n654), .Y (y79) );
  OAI21xp33_ASAP7_75t_R  g392( .A1 (n654), .A2 (n655), .B (n657), .Y (n660) );
  NOR2xp33_ASAP7_75t_R   g393( .A (x80), .B (x208), .Y (n661) );
  AND2x2_ASAP7_75t_R     g394( .A (x80), .B (x208), .Y (n662) );
  NOR2xp33_ASAP7_75t_R   g395( .A (n661), .B (n662), .Y (n663) );
  XOR2xp5_ASAP7_75t_R    g396( .A (n660), .B (n663), .Y (y80) );
  MAJIxp5_ASAP7_75t_R    g397( .A (n660), .B (x208), .C (x80), .Y (n665) );
  NOR2xp33_ASAP7_75t_R   g398( .A (x81), .B (x209), .Y (n666) );
  NAND2xp33_ASAP7_75t_R  g399( .A (x81), .B (x209), .Y (n667) );
  INVx1_ASAP7_75t_R      g400( .A (n667), .Y (n668) );
  NOR2xp33_ASAP7_75t_R   g401( .A (n666), .B (n668), .Y (n669) );
  XNOR2xp5_ASAP7_75t_R   g402( .A (n665), .B (n669), .Y (y81) );
  OAI21xp33_ASAP7_75t_R  g403( .A1 (n665), .A2 (n666), .B (n667), .Y (n671) );
  NOR2xp33_ASAP7_75t_R   g404( .A (x82), .B (x210), .Y (n672) );
  AND2x2_ASAP7_75t_R     g405( .A (x82), .B (x210), .Y (n673) );
  NOR2xp33_ASAP7_75t_R   g406( .A (n672), .B (n673), .Y (n674) );
  XOR2xp5_ASAP7_75t_R    g407( .A (n671), .B (n674), .Y (y82) );
  MAJIxp5_ASAP7_75t_R    g408( .A (n671), .B (x210), .C (x82), .Y (n676) );
  NOR2xp33_ASAP7_75t_R   g409( .A (x83), .B (x211), .Y (n677) );
  NAND2xp33_ASAP7_75t_R  g410( .A (x83), .B (x211), .Y (n678) );
  INVx1_ASAP7_75t_R      g411( .A (n678), .Y (n679) );
  NOR2xp33_ASAP7_75t_R   g412( .A (n677), .B (n679), .Y (n680) );
  XNOR2xp5_ASAP7_75t_R   g413( .A (n676), .B (n680), .Y (y83) );
  OAI21xp33_ASAP7_75t_R  g414( .A1 (n676), .A2 (n677), .B (n678), .Y (n682) );
  NOR2xp33_ASAP7_75t_R   g415( .A (x84), .B (x212), .Y (n683) );
  AND2x2_ASAP7_75t_R     g416( .A (x84), .B (x212), .Y (n684) );
  NOR2xp33_ASAP7_75t_R   g417( .A (n683), .B (n684), .Y (n685) );
  XOR2xp5_ASAP7_75t_R    g418( .A (n682), .B (n685), .Y (y84) );
  MAJIxp5_ASAP7_75t_R    g419( .A (n682), .B (x212), .C (x84), .Y (n687) );
  XOR2xp5_ASAP7_75t_R    g420( .A (x85), .B (x213), .Y (n688) );
  XNOR2xp5_ASAP7_75t_R   g421( .A (n687), .B (n688), .Y (y85) );
  INVx1_ASAP7_75t_R      g422( .A (x85), .Y (n264) );
  INVx1_ASAP7_75t_R      g423( .A (x213), .Y (n275) );
  MAJIxp5_ASAP7_75t_R    g424( .A (n264), .B (n275), .C (n687), .Y (n690) );
  NOR2xp33_ASAP7_75t_R   g425( .A (x86), .B (x214), .Y (n691) );
  AND2x2_ASAP7_75t_R     g426( .A (x86), .B (x214), .Y (n692) );
  NOR2xp33_ASAP7_75t_R   g427( .A (n691), .B (n692), .Y (n693) );
  XOR2xp5_ASAP7_75t_R    g428( .A (n690), .B (n693), .Y (y86) );
  NOR2xp33_ASAP7_75t_R   g429( .A (x87), .B (x215), .Y (n696) );
  INVx1_ASAP7_75t_R      g430( .A (n696), .Y (n697) );
  NAND2xp33_ASAP7_75t_R  g431( .A (x87), .B (x215), .Y (n698) );
  NAND2xp33_ASAP7_75t_R  g432( .A (n697), .B (n698), .Y (n699) );
  MAJIxp5_ASAP7_75t_R    g433( .A (n690), .B (x214), .C (x86), .Y (n695) );
  XOR2xp5_ASAP7_75t_R    g434( .A (n699), .B (n695), .Y (y87) );
  OAI21xp33_ASAP7_75t_R  g435( .A1 (n695), .A2 (n696), .B (n698), .Y (n701) );
  XOR2xp5_ASAP7_75t_R    g436( .A (x88), .B (x216), .Y (n702) );
  XOR2xp5_ASAP7_75t_R    g437( .A (n701), .B (n702), .Y (y88) );
  MAJIxp5_ASAP7_75t_R    g438( .A (n701), .B (x216), .C (x88), .Y (n704) );
  NOR2xp33_ASAP7_75t_R   g439( .A (x89), .B (x217), .Y (n705) );
  NAND2xp33_ASAP7_75t_R  g440( .A (x89), .B (x217), .Y (n706) );
  INVx1_ASAP7_75t_R      g441( .A (n706), .Y (n707) );
  NOR2xp33_ASAP7_75t_R   g442( .A (n705), .B (n707), .Y (n708) );
  XNOR2xp5_ASAP7_75t_R   g443( .A (n704), .B (n708), .Y (y89) );
  OAI21xp33_ASAP7_75t_R  g444( .A1 (n704), .A2 (n705), .B (n706), .Y (n710) );
  XOR2xp5_ASAP7_75t_R    g445( .A (x90), .B (x218), .Y (n711) );
  XOR2xp5_ASAP7_75t_R    g446( .A (n710), .B (n711), .Y (y90) );
  MAJIxp5_ASAP7_75t_R    g447( .A (n710), .B (x218), .C (x90), .Y (n713) );
  NOR2xp33_ASAP7_75t_R   g448( .A (x91), .B (x219), .Y (n714) );
  NAND2xp33_ASAP7_75t_R  g449( .A (x91), .B (x219), .Y (n715) );
  INVx1_ASAP7_75t_R      g450( .A (n715), .Y (n716) );
  NOR2xp33_ASAP7_75t_R   g451( .A (n714), .B (n716), .Y (n717) );
  XNOR2xp5_ASAP7_75t_R   g452( .A (n713), .B (n717), .Y (y91) );
  OAI21xp33_ASAP7_75t_R  g453( .A1 (n713), .A2 (n714), .B (n715), .Y (n719) );
  XOR2xp5_ASAP7_75t_R    g454( .A (x92), .B (x220), .Y (n720) );
  XOR2xp5_ASAP7_75t_R    g455( .A (n719), .B (n720), .Y (y92) );
  MAJIxp5_ASAP7_75t_R    g456( .A (n719), .B (x220), .C (x92), .Y (n722) );
  NOR2xp33_ASAP7_75t_R   g457( .A (x93), .B (x221), .Y (n723) );
  NAND2xp33_ASAP7_75t_R  g458( .A (x93), .B (x221), .Y (n724) );
  INVx1_ASAP7_75t_R      g459( .A (n724), .Y (n725) );
  NOR2xp33_ASAP7_75t_R   g460( .A (n723), .B (n725), .Y (n726) );
  XNOR2xp5_ASAP7_75t_R   g461( .A (n722), .B (n726), .Y (y93) );
  OAI21xp33_ASAP7_75t_R  g462( .A1 (n722), .A2 (n723), .B (n724), .Y (n728) );
  XNOR2xp5_ASAP7_75t_R   g463( .A (x94), .B (x222), .Y (n729) );
  XNOR2xp5_ASAP7_75t_R   g464( .A (n728), .B (n729), .Y (y94) );
  NOR2xp33_ASAP7_75t_R   g465( .A (x95), .B (x223), .Y (n732) );
  INVx1_ASAP7_75t_R      g466( .A (n732), .Y (n733) );
  NAND2xp33_ASAP7_75t_R  g467( .A (x95), .B (x223), .Y (n734) );
  NAND2xp33_ASAP7_75t_R  g468( .A (n733), .B (n734), .Y (n735) );
  MAJIxp5_ASAP7_75t_R    g469( .A (n728), .B (x222), .C (x94), .Y (n731) );
  XOR2xp5_ASAP7_75t_R    g470( .A (n735), .B (n731), .Y (y95) );
  OAI21xp33_ASAP7_75t_R  g471( .A1 (n731), .A2 (n732), .B (n734), .Y (n737) );
  NOR2xp33_ASAP7_75t_R   g472( .A (x96), .B (x224), .Y (n738) );
  AND2x2_ASAP7_75t_R     g473( .A (x96), .B (x224), .Y (n739) );
  NOR2xp33_ASAP7_75t_R   g474( .A (n738), .B (n739), .Y (n740) );
  XOR2xp5_ASAP7_75t_R    g475( .A (n737), .B (n740), .Y (y96) );
  MAJIxp5_ASAP7_75t_R    g476( .A (n737), .B (x224), .C (x96), .Y (n742) );
  NOR2xp33_ASAP7_75t_R   g477( .A (x97), .B (x225), .Y (n743) );
  NAND2xp33_ASAP7_75t_R  g478( .A (x97), .B (x225), .Y (n744) );
  INVx1_ASAP7_75t_R      g479( .A (n744), .Y (n745) );
  NOR2xp33_ASAP7_75t_R   g480( .A (n743), .B (n745), .Y (n746) );
  XNOR2xp5_ASAP7_75t_R   g481( .A (n742), .B (n746), .Y (y97) );
  OAI21xp33_ASAP7_75t_R  g482( .A1 (n742), .A2 (n743), .B (n744), .Y (n748) );
  XOR2xp5_ASAP7_75t_R    g483( .A (x98), .B (x226), .Y (n749) );
  XOR2xp5_ASAP7_75t_R    g484( .A (n748), .B (n749), .Y (y98) );
  MAJIxp5_ASAP7_75t_R    g485( .A (n748), .B (x226), .C (x98), .Y (n751) );
  NOR2xp33_ASAP7_75t_R   g486( .A (x99), .B (x227), .Y (n752) );
  NAND2xp33_ASAP7_75t_R  g487( .A (x99), .B (x227), .Y (n753) );
  INVx1_ASAP7_75t_R      g488( .A (n753), .Y (n754) );
  NOR2xp33_ASAP7_75t_R   g489( .A (n752), .B (n754), .Y (n755) );
  XNOR2xp5_ASAP7_75t_R   g490( .A (n751), .B (n755), .Y (y99) );
  OAI21xp33_ASAP7_75t_R  g491( .A1 (n751), .A2 (n752), .B (n753), .Y (n757) );
  XNOR2xp5_ASAP7_75t_R   g492( .A (x100), .B (x228), .Y (n758) );
  XNOR2xp5_ASAP7_75t_R   g493( .A (n757), .B (n758), .Y (y100) );
  NOR2xp33_ASAP7_75t_R   g494( .A (x101), .B (x229), .Y (n761) );
  INVx1_ASAP7_75t_R      g495( .A (n761), .Y (n762) );
  NAND2xp33_ASAP7_75t_R  g496( .A (x101), .B (x229), .Y (n763) );
  NAND2xp33_ASAP7_75t_R  g497( .A (n762), .B (n763), .Y (n764) );
  MAJIxp5_ASAP7_75t_R    g498( .A (n757), .B (x228), .C (x100), .Y (n760) );
  XOR2xp5_ASAP7_75t_R    g499( .A (n764), .B (n760), .Y (y101) );
  OAI21xp33_ASAP7_75t_R  g500( .A1 (n760), .A2 (n761), .B (n763), .Y (n766) );
  NOR2xp33_ASAP7_75t_R   g501( .A (x102), .B (x230), .Y (n767) );
  AND2x2_ASAP7_75t_R     g502( .A (x102), .B (x230), .Y (n768) );
  NOR2xp33_ASAP7_75t_R   g503( .A (n767), .B (n768), .Y (n769) );
  XOR2xp5_ASAP7_75t_R    g504( .A (n766), .B (n769), .Y (y102) );
  MAJIxp5_ASAP7_75t_R    g505( .A (n766), .B (x230), .C (x102), .Y (n771) );
  XOR2xp5_ASAP7_75t_R    g506( .A (x103), .B (x231), .Y (n772) );
  XNOR2xp5_ASAP7_75t_R   g507( .A (n771), .B (n772), .Y (y103) );
  INVx1_ASAP7_75t_R      g508( .A (x103), .Y (n265) );
  INVx1_ASAP7_75t_R      g509( .A (x231), .Y (n276) );
  MAJIxp5_ASAP7_75t_R    g510( .A (n265), .B (n276), .C (n771), .Y (n774) );
  XOR2xp5_ASAP7_75t_R    g511( .A (x104), .B (x232), .Y (n775) );
  XOR2xp5_ASAP7_75t_R    g512( .A (n774), .B (n775), .Y (y104) );
  NOR2xp33_ASAP7_75t_R   g513( .A (x105), .B (x233), .Y (n778) );
  INVx1_ASAP7_75t_R      g514( .A (n778), .Y (n779) );
  NAND2xp33_ASAP7_75t_R  g515( .A (x105), .B (x233), .Y (n780) );
  NAND2xp33_ASAP7_75t_R  g516( .A (n779), .B (n780), .Y (n781) );
  MAJIxp5_ASAP7_75t_R    g517( .A (n774), .B (x232), .C (x104), .Y (n777) );
  XOR2xp5_ASAP7_75t_R    g518( .A (n781), .B (n777), .Y (y105) );
  OAI21xp33_ASAP7_75t_R  g519( .A1 (n777), .A2 (n778), .B (n780), .Y (n783) );
  NOR2xp33_ASAP7_75t_R   g520( .A (x106), .B (x234), .Y (n784) );
  AND2x2_ASAP7_75t_R     g521( .A (x106), .B (x234), .Y (n785) );
  NOR2xp33_ASAP7_75t_R   g522( .A (n784), .B (n785), .Y (n786) );
  XOR2xp5_ASAP7_75t_R    g523( .A (n783), .B (n786), .Y (y106) );
  MAJIxp5_ASAP7_75t_R    g524( .A (n783), .B (x234), .C (x106), .Y (n788) );
  XOR2xp5_ASAP7_75t_R    g525( .A (x107), .B (x235), .Y (n789) );
  XNOR2xp5_ASAP7_75t_R   g526( .A (n788), .B (n789), .Y (y107) );
  INVx1_ASAP7_75t_R      g527( .A (x107), .Y (n266) );
  INVx1_ASAP7_75t_R      g528( .A (x235), .Y (n277) );
  MAJIxp5_ASAP7_75t_R    g529( .A (n266), .B (n277), .C (n788), .Y (n791) );
  OR2x2_ASAP7_75t_R      g530( .A (x108), .B (x236), .Y (n792) );
  NAND2xp33_ASAP7_75t_R  g531( .A (x108), .B (x236), .Y (n793) );
  NAND2xp33_ASAP7_75t_R  g532( .A (n792), .B (n793), .Y (n794) );
  XNOR2xp5_ASAP7_75t_R   g533( .A (n791), .B (n794), .Y (y108) );
  NOR2xp33_ASAP7_75t_R   g534( .A (x109), .B (x237), .Y (n797) );
  INVx1_ASAP7_75t_R      g535( .A (n797), .Y (n798) );
  NAND2xp33_ASAP7_75t_R  g536( .A (x109), .B (x237), .Y (n799) );
  NAND2xp33_ASAP7_75t_R  g537( .A (n798), .B (n799), .Y (n800) );
  MAJIxp5_ASAP7_75t_R    g538( .A (n791), .B (x236), .C (x108), .Y (n796) );
  XOR2xp5_ASAP7_75t_R    g539( .A (n800), .B (n796), .Y (y109) );
  OAI21xp33_ASAP7_75t_R  g540( .A1 (n796), .A2 (n797), .B (n799), .Y (n802) );
  XNOR2xp5_ASAP7_75t_R   g541( .A (x110), .B (x238), .Y (n803) );
  XNOR2xp5_ASAP7_75t_R   g542( .A (n802), .B (n803), .Y (y110) );
  MAJIxp5_ASAP7_75t_R    g543( .A (n802), .B (x238), .C (x110), .Y (n805) );
  NOR2xp33_ASAP7_75t_R   g544( .A (x111), .B (x239), .Y (n806) );
  NAND2xp33_ASAP7_75t_R  g545( .A (x111), .B (x239), .Y (n807) );
  INVx1_ASAP7_75t_R      g546( .A (n807), .Y (n808) );
  NOR2xp33_ASAP7_75t_R   g547( .A (n806), .B (n808), .Y (n809) );
  XNOR2xp5_ASAP7_75t_R   g548( .A (n805), .B (n809), .Y (y111) );
  OAI21xp33_ASAP7_75t_R  g549( .A1 (n805), .A2 (n806), .B (n807), .Y (n811) );
  NOR2xp33_ASAP7_75t_R   g550( .A (x112), .B (x240), .Y (n812) );
  AND2x2_ASAP7_75t_R     g551( .A (x112), .B (x240), .Y (n813) );
  NOR2xp33_ASAP7_75t_R   g552( .A (n812), .B (n813), .Y (n814) );
  XOR2xp5_ASAP7_75t_R    g553( .A (n811), .B (n814), .Y (y112) );
  MAJIxp5_ASAP7_75t_R    g554( .A (n811), .B (x240), .C (x112), .Y (n816) );
  XOR2xp5_ASAP7_75t_R    g555( .A (x113), .B (x241), .Y (n817) );
  XNOR2xp5_ASAP7_75t_R   g556( .A (n816), .B (n817), .Y (y113) );
  INVx1_ASAP7_75t_R      g557( .A (x113), .Y (n267) );
  INVx1_ASAP7_75t_R      g558( .A (x241), .Y (n278) );
  MAJIxp5_ASAP7_75t_R    g559( .A (n267), .B (n278), .C (n816), .Y (n819) );
  XNOR2xp5_ASAP7_75t_R   g560( .A (x114), .B (x242), .Y (n820) );
  XNOR2xp5_ASAP7_75t_R   g561( .A (n819), .B (n820), .Y (y114) );
  NOR2xp33_ASAP7_75t_R   g562( .A (x115), .B (x243), .Y (n823) );
  INVx1_ASAP7_75t_R      g563( .A (n823), .Y (n824) );
  NAND2xp33_ASAP7_75t_R  g564( .A (x115), .B (x243), .Y (n825) );
  NAND2xp33_ASAP7_75t_R  g565( .A (n824), .B (n825), .Y (n826) );
  MAJIxp5_ASAP7_75t_R    g566( .A (n819), .B (x242), .C (x114), .Y (n822) );
  XOR2xp5_ASAP7_75t_R    g567( .A (n826), .B (n822), .Y (y115) );
  OAI21xp33_ASAP7_75t_R  g568( .A1 (n822), .A2 (n823), .B (n825), .Y (n828) );
  NOR2xp33_ASAP7_75t_R   g569( .A (x116), .B (x244), .Y (n829) );
  AND2x2_ASAP7_75t_R     g570( .A (x116), .B (x244), .Y (n830) );
  NOR2xp33_ASAP7_75t_R   g571( .A (n829), .B (n830), .Y (n831) );
  XOR2xp5_ASAP7_75t_R    g572( .A (n828), .B (n831), .Y (y116) );
  MAJIxp5_ASAP7_75t_R    g573( .A (n828), .B (x244), .C (x116), .Y (n833) );
  NOR2xp33_ASAP7_75t_R   g574( .A (x117), .B (x245), .Y (n834) );
  NAND2xp33_ASAP7_75t_R  g575( .A (x117), .B (x245), .Y (n835) );
  INVx1_ASAP7_75t_R      g576( .A (n835), .Y (n836) );
  NOR2xp33_ASAP7_75t_R   g577( .A (n834), .B (n836), .Y (n837) );
  XNOR2xp5_ASAP7_75t_R   g578( .A (n833), .B (n837), .Y (y117) );
  OAI21xp33_ASAP7_75t_R  g579( .A1 (n833), .A2 (n834), .B (n835), .Y (n839) );
  NOR2xp33_ASAP7_75t_R   g580( .A (x118), .B (x246), .Y (n840) );
  AND2x2_ASAP7_75t_R     g581( .A (x118), .B (x246), .Y (n841) );
  NOR2xp33_ASAP7_75t_R   g582( .A (n840), .B (n841), .Y (n842) );
  XOR2xp5_ASAP7_75t_R    g583( .A (n839), .B (n842), .Y (y118) );
  MAJIxp5_ASAP7_75t_R    g584( .A (n839), .B (x246), .C (x118), .Y (n844) );
  NOR2xp33_ASAP7_75t_R   g585( .A (x119), .B (x247), .Y (n845) );
  NAND2xp33_ASAP7_75t_R  g586( .A (x119), .B (x247), .Y (n846) );
  INVx1_ASAP7_75t_R      g587( .A (n846), .Y (n847) );
  NOR2xp33_ASAP7_75t_R   g588( .A (n845), .B (n847), .Y (n848) );
  XNOR2xp5_ASAP7_75t_R   g589( .A (n844), .B (n848), .Y (y119) );
  OAI21xp33_ASAP7_75t_R  g590( .A1 (n844), .A2 (n845), .B (n846), .Y (n850) );
  NOR2xp33_ASAP7_75t_R   g591( .A (x120), .B (x248), .Y (n851) );
  AND2x2_ASAP7_75t_R     g592( .A (x120), .B (x248), .Y (n852) );
  NOR2xp33_ASAP7_75t_R   g593( .A (n851), .B (n852), .Y (n853) );
  XOR2xp5_ASAP7_75t_R    g594( .A (n850), .B (n853), .Y (y120) );
  MAJIxp5_ASAP7_75t_R    g595( .A (n850), .B (x248), .C (x120), .Y (n855) );
  NOR2xp33_ASAP7_75t_R   g596( .A (x121), .B (x249), .Y (n856) );
  NAND2xp33_ASAP7_75t_R  g597( .A (x121), .B (x249), .Y (n857) );
  INVx1_ASAP7_75t_R      g598( .A (n857), .Y (n858) );
  NOR2xp33_ASAP7_75t_R   g599( .A (n856), .B (n858), .Y (n859) );
  XNOR2xp5_ASAP7_75t_R   g600( .A (n855), .B (n859), .Y (y121) );
  OAI21xp33_ASAP7_75t_R  g601( .A1 (n855), .A2 (n856), .B (n857), .Y (n861) );
  NOR2xp33_ASAP7_75t_R   g602( .A (x122), .B (x250), .Y (n862) );
  AND2x2_ASAP7_75t_R     g603( .A (x122), .B (x250), .Y (n863) );
  NOR2xp33_ASAP7_75t_R   g604( .A (n862), .B (n863), .Y (n864) );
  XOR2xp5_ASAP7_75t_R    g605( .A (n861), .B (n864), .Y (y122) );
  MAJIxp5_ASAP7_75t_R    g606( .A (n861), .B (x250), .C (x122), .Y (n866) );
  NOR2xp33_ASAP7_75t_R   g607( .A (x123), .B (x251), .Y (n867) );
  NAND2xp33_ASAP7_75t_R  g608( .A (x123), .B (x251), .Y (n868) );
  INVx1_ASAP7_75t_R      g609( .A (n868), .Y (n869) );
  NOR2xp33_ASAP7_75t_R   g610( .A (n867), .B (n869), .Y (n870) );
  XNOR2xp5_ASAP7_75t_R   g611( .A (n866), .B (n870), .Y (y123) );
  OAI21xp33_ASAP7_75t_R  g612( .A1 (n866), .A2 (n867), .B (n868), .Y (n872) );
  XOR2xp5_ASAP7_75t_R    g613( .A (x124), .B (x252), .Y (n873) );
  XOR2xp5_ASAP7_75t_R    g614( .A (n872), .B (n873), .Y (y124) );
  MAJIxp5_ASAP7_75t_R    g615( .A (n872), .B (x252), .C (x124), .Y (n875) );
  XOR2xp5_ASAP7_75t_R    g616( .A (x125), .B (x253), .Y (n876) );
  XNOR2xp5_ASAP7_75t_R   g617( .A (n875), .B (n876), .Y (y125) );
  INVx1_ASAP7_75t_R      g618( .A (x125), .Y (n268) );
  INVx1_ASAP7_75t_R      g619( .A (x253), .Y (n279) );
  MAJIxp5_ASAP7_75t_R    g620( .A (n268), .B (n279), .C (n875), .Y (n878) );
  NOR2xp33_ASAP7_75t_R   g621( .A (x126), .B (x254), .Y (n879) );
  AND2x2_ASAP7_75t_R     g622( .A (x126), .B (x254), .Y (n880) );
  NOR2xp33_ASAP7_75t_R   g623( .A (n879), .B (n880), .Y (n881) );
  XOR2xp5_ASAP7_75t_R    g624( .A (n878), .B (n881), .Y (y126) );
  MAJIxp5_ASAP7_75t_R    g625( .A (n878), .B (x254), .C (x126), .Y (n883) );
  NOR2xp33_ASAP7_75t_R   g626( .A (x127), .B (x255), .Y (n884) );
  NAND2xp33_ASAP7_75t_R  g627( .A (x127), .B (x255), .Y (n885) );
  INVx1_ASAP7_75t_R      g628( .A (n885), .Y (n886) );
  NOR2xp33_ASAP7_75t_R   g629( .A (n884), .B (n886), .Y (n887) );
  XNOR2xp5_ASAP7_75t_R   g630( .A (n883), .B (n887), .Y (y127) );
  OAI21xp33_ASAP7_75t_R  g631( .A1 (n883), .A2 (n884), .B (n885), .Y (y128) );
endmodule
