module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 ;
  wire n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n515 , n516 , n517 , n518 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1643 , n1644 , n1645 , n1646 , n1647 , n1649 ;
  INVx1_ASAP7_75t_R      g0000( .A (x0), .Y (n258) );
  XNOR2xp5_ASAP7_75t_R   g0001( .A (n258), .B (x128), .Y (y0) );
  NAND2xp33_ASAP7_75t_R  g0002( .A (x0), .B (x128), .Y (n515) );
  INVx1_ASAP7_75t_R      g0003( .A (x1), .Y (n259) );
  XNOR2xp5_ASAP7_75t_R   g0004( .A (n259), .B (x129), .Y (n518) );
  XNOR2xp5_ASAP7_75t_R   g0005( .A (n515), .B (n518), .Y (y1) );
  INVx1_ASAP7_75t_R      g0006( .A (x129), .Y (n387) );
  NOR2xp33_ASAP7_75t_R   g0007( .A (n259), .B (n387), .Y (n516) );
  INVx1_ASAP7_75t_R      g0008( .A (x128), .Y (n386) );
  AOI211xp5_ASAP7_75t_R  g0009( .A1 (n259), .B (n386), .C (n258), .A2 (n387), .Y (n520) );
  NOR2xp33_ASAP7_75t_R   g0010( .A (n516), .B (n520), .Y (n522) );
  INVx1_ASAP7_75t_R      g0011( .A (x2), .Y (n260) );
  XNOR2xp5_ASAP7_75t_R   g0012( .A (n260), .B (x130), .Y (n527) );
  XNOR2xp5_ASAP7_75t_R   g0013( .A (n522), .B (n527), .Y (y2) );
  INVx1_ASAP7_75t_R      g0014( .A (x130), .Y (n388) );
  NOR2xp33_ASAP7_75t_R   g0015( .A (n260), .B (n388), .Y (n525) );
  NAND2xp33_ASAP7_75t_R  g0016( .A (x1), .B (x129), .Y (n517) );
  NOR2xp33_ASAP7_75t_R   g0017( .A (x2), .B (x130), .Y (n523) );
  OAI211xp5_ASAP7_75t_R  g0018( .A1 (x1), .A2 (x129), .B (x128), .C (x0), .Y (n521) );
  AOI21xp33_ASAP7_75t_R  g0019( .A1 (n517), .B (n523), .A2 (n521), .Y (n529) );
  NOR2xp33_ASAP7_75t_R   g0020( .A (n525), .B (n529), .Y (n531) );
  INVx1_ASAP7_75t_R      g0021( .A (x3), .Y (n261) );
  XNOR2xp5_ASAP7_75t_R   g0022( .A (n261), .B (x131), .Y (n536) );
  XNOR2xp5_ASAP7_75t_R   g0023( .A (n531), .B (n536), .Y (y3) );
  INVx1_ASAP7_75t_R      g0024( .A (x131), .Y (n389) );
  NOR2xp33_ASAP7_75t_R   g0025( .A (n261), .B (n389), .Y (n534) );
  NAND2xp33_ASAP7_75t_R  g0026( .A (x2), .B (x130), .Y (n526) );
  NOR2xp33_ASAP7_75t_R   g0027( .A (x3), .B (x131), .Y (n532) );
  NAND2xp33_ASAP7_75t_R  g0028( .A (n260), .B (n388), .Y (n524) );
  OAI21xp33_ASAP7_75t_R  g0029( .A1 (n516), .A2 (n520), .B (n524), .Y (n530) );
  AOI21xp33_ASAP7_75t_R  g0030( .A1 (n526), .B (n532), .A2 (n530), .Y (n538) );
  NOR2xp33_ASAP7_75t_R   g0031( .A (n534), .B (n538), .Y (n540) );
  INVx1_ASAP7_75t_R      g0032( .A (x4), .Y (n262) );
  XNOR2xp5_ASAP7_75t_R   g0033( .A (n262), .B (x132), .Y (n545) );
  XNOR2xp5_ASAP7_75t_R   g0034( .A (n540), .B (n545), .Y (y4) );
  INVx1_ASAP7_75t_R      g0035( .A (x132), .Y (n390) );
  NOR2xp33_ASAP7_75t_R   g0036( .A (n262), .B (n390), .Y (n543) );
  NAND2xp33_ASAP7_75t_R  g0037( .A (x3), .B (x131), .Y (n535) );
  NOR2xp33_ASAP7_75t_R   g0038( .A (x4), .B (x132), .Y (n541) );
  NAND2xp33_ASAP7_75t_R  g0039( .A (n261), .B (n389), .Y (n533) );
  OAI21xp33_ASAP7_75t_R  g0040( .A1 (n525), .A2 (n529), .B (n533), .Y (n539) );
  AOI21xp33_ASAP7_75t_R  g0041( .A1 (n535), .B (n541), .A2 (n539), .Y (n547) );
  NOR2xp33_ASAP7_75t_R   g0042( .A (n543), .B (n547), .Y (n549) );
  INVx1_ASAP7_75t_R      g0043( .A (x5), .Y (n263) );
  XNOR2xp5_ASAP7_75t_R   g0044( .A (n263), .B (x133), .Y (n554) );
  XNOR2xp5_ASAP7_75t_R   g0045( .A (n549), .B (n554), .Y (y5) );
  INVx1_ASAP7_75t_R      g0046( .A (x133), .Y (n391) );
  NOR2xp33_ASAP7_75t_R   g0047( .A (n263), .B (n391), .Y (n552) );
  NAND2xp33_ASAP7_75t_R  g0048( .A (x4), .B (x132), .Y (n544) );
  NOR2xp33_ASAP7_75t_R   g0049( .A (x5), .B (x133), .Y (n550) );
  NAND2xp33_ASAP7_75t_R  g0050( .A (n262), .B (n390), .Y (n542) );
  OAI21xp33_ASAP7_75t_R  g0051( .A1 (n534), .A2 (n538), .B (n542), .Y (n548) );
  AOI21xp33_ASAP7_75t_R  g0052( .A1 (n544), .B (n550), .A2 (n548), .Y (n556) );
  NOR2xp33_ASAP7_75t_R   g0053( .A (n552), .B (n556), .Y (n558) );
  INVx1_ASAP7_75t_R      g0054( .A (x6), .Y (n264) );
  XNOR2xp5_ASAP7_75t_R   g0055( .A (n264), .B (x134), .Y (n563) );
  XNOR2xp5_ASAP7_75t_R   g0056( .A (n558), .B (n563), .Y (y6) );
  INVx1_ASAP7_75t_R      g0057( .A (x134), .Y (n392) );
  NOR2xp33_ASAP7_75t_R   g0058( .A (n264), .B (n392), .Y (n561) );
  NAND2xp33_ASAP7_75t_R  g0059( .A (x5), .B (x133), .Y (n553) );
  NOR2xp33_ASAP7_75t_R   g0060( .A (x6), .B (x134), .Y (n559) );
  NAND2xp33_ASAP7_75t_R  g0061( .A (n263), .B (n391), .Y (n551) );
  OAI21xp33_ASAP7_75t_R  g0062( .A1 (n543), .A2 (n547), .B (n551), .Y (n557) );
  AOI21xp33_ASAP7_75t_R  g0063( .A1 (n553), .B (n559), .A2 (n557), .Y (n565) );
  NOR2xp33_ASAP7_75t_R   g0064( .A (n561), .B (n565), .Y (n567) );
  INVx1_ASAP7_75t_R      g0065( .A (x7), .Y (n265) );
  XNOR2xp5_ASAP7_75t_R   g0066( .A (n265), .B (x135), .Y (n572) );
  XNOR2xp5_ASAP7_75t_R   g0067( .A (n567), .B (n572), .Y (y7) );
  INVx1_ASAP7_75t_R      g0068( .A (x135), .Y (n393) );
  NOR2xp33_ASAP7_75t_R   g0069( .A (n265), .B (n393), .Y (n570) );
  NAND2xp33_ASAP7_75t_R  g0070( .A (x6), .B (x134), .Y (n562) );
  NOR2xp33_ASAP7_75t_R   g0071( .A (x7), .B (x135), .Y (n568) );
  NAND2xp33_ASAP7_75t_R  g0072( .A (n264), .B (n392), .Y (n560) );
  OAI21xp33_ASAP7_75t_R  g0073( .A1 (n552), .A2 (n556), .B (n560), .Y (n566) );
  AOI21xp33_ASAP7_75t_R  g0074( .A1 (n562), .B (n568), .A2 (n566), .Y (n574) );
  NOR2xp33_ASAP7_75t_R   g0075( .A (n570), .B (n574), .Y (n576) );
  INVx1_ASAP7_75t_R      g0076( .A (x8), .Y (n266) );
  XNOR2xp5_ASAP7_75t_R   g0077( .A (n266), .B (x136), .Y (n581) );
  XNOR2xp5_ASAP7_75t_R   g0078( .A (n576), .B (n581), .Y (y8) );
  INVx1_ASAP7_75t_R      g0079( .A (x136), .Y (n394) );
  NOR2xp33_ASAP7_75t_R   g0080( .A (n266), .B (n394), .Y (n579) );
  NAND2xp33_ASAP7_75t_R  g0081( .A (x7), .B (x135), .Y (n571) );
  NOR2xp33_ASAP7_75t_R   g0082( .A (x8), .B (x136), .Y (n577) );
  NAND2xp33_ASAP7_75t_R  g0083( .A (n265), .B (n393), .Y (n569) );
  OAI21xp33_ASAP7_75t_R  g0084( .A1 (n561), .A2 (n565), .B (n569), .Y (n575) );
  AOI21xp33_ASAP7_75t_R  g0085( .A1 (n571), .B (n577), .A2 (n575), .Y (n583) );
  NOR2xp33_ASAP7_75t_R   g0086( .A (n579), .B (n583), .Y (n585) );
  INVx1_ASAP7_75t_R      g0087( .A (x9), .Y (n267) );
  XNOR2xp5_ASAP7_75t_R   g0088( .A (n267), .B (x137), .Y (n590) );
  XNOR2xp5_ASAP7_75t_R   g0089( .A (n585), .B (n590), .Y (y9) );
  INVx1_ASAP7_75t_R      g0090( .A (x137), .Y (n395) );
  NOR2xp33_ASAP7_75t_R   g0091( .A (n267), .B (n395), .Y (n588) );
  NAND2xp33_ASAP7_75t_R  g0092( .A (x8), .B (x136), .Y (n580) );
  NOR2xp33_ASAP7_75t_R   g0093( .A (x9), .B (x137), .Y (n586) );
  NAND2xp33_ASAP7_75t_R  g0094( .A (n266), .B (n394), .Y (n578) );
  OAI21xp33_ASAP7_75t_R  g0095( .A1 (n570), .A2 (n574), .B (n578), .Y (n584) );
  AOI21xp33_ASAP7_75t_R  g0096( .A1 (n580), .B (n586), .A2 (n584), .Y (n592) );
  NOR2xp33_ASAP7_75t_R   g0097( .A (n588), .B (n592), .Y (n594) );
  INVx1_ASAP7_75t_R      g0098( .A (x10), .Y (n268) );
  XNOR2xp5_ASAP7_75t_R   g0099( .A (n268), .B (x138), .Y (n599) );
  XNOR2xp5_ASAP7_75t_R   g0100( .A (n594), .B (n599), .Y (y10) );
  INVx1_ASAP7_75t_R      g0101( .A (x138), .Y (n396) );
  NOR2xp33_ASAP7_75t_R   g0102( .A (n268), .B (n396), .Y (n597) );
  NAND2xp33_ASAP7_75t_R  g0103( .A (x9), .B (x137), .Y (n589) );
  NOR2xp33_ASAP7_75t_R   g0104( .A (x10), .B (x138), .Y (n595) );
  NAND2xp33_ASAP7_75t_R  g0105( .A (n267), .B (n395), .Y (n587) );
  OAI21xp33_ASAP7_75t_R  g0106( .A1 (n579), .A2 (n583), .B (n587), .Y (n593) );
  AOI21xp33_ASAP7_75t_R  g0107( .A1 (n589), .B (n595), .A2 (n593), .Y (n601) );
  NOR2xp33_ASAP7_75t_R   g0108( .A (n597), .B (n601), .Y (n603) );
  INVx1_ASAP7_75t_R      g0109( .A (x11), .Y (n269) );
  XNOR2xp5_ASAP7_75t_R   g0110( .A (n269), .B (x139), .Y (n608) );
  XNOR2xp5_ASAP7_75t_R   g0111( .A (n603), .B (n608), .Y (y11) );
  INVx1_ASAP7_75t_R      g0112( .A (x139), .Y (n397) );
  NOR2xp33_ASAP7_75t_R   g0113( .A (n269), .B (n397), .Y (n606) );
  NAND2xp33_ASAP7_75t_R  g0114( .A (x10), .B (x138), .Y (n598) );
  NOR2xp33_ASAP7_75t_R   g0115( .A (x11), .B (x139), .Y (n604) );
  NAND2xp33_ASAP7_75t_R  g0116( .A (n268), .B (n396), .Y (n596) );
  OAI21xp33_ASAP7_75t_R  g0117( .A1 (n588), .A2 (n592), .B (n596), .Y (n602) );
  AOI21xp33_ASAP7_75t_R  g0118( .A1 (n598), .B (n604), .A2 (n602), .Y (n610) );
  NOR2xp33_ASAP7_75t_R   g0119( .A (n606), .B (n610), .Y (n612) );
  INVx1_ASAP7_75t_R      g0120( .A (x12), .Y (n270) );
  XNOR2xp5_ASAP7_75t_R   g0121( .A (n270), .B (x140), .Y (n617) );
  XNOR2xp5_ASAP7_75t_R   g0122( .A (n612), .B (n617), .Y (y12) );
  INVx1_ASAP7_75t_R      g0123( .A (x140), .Y (n398) );
  NOR2xp33_ASAP7_75t_R   g0124( .A (n270), .B (n398), .Y (n615) );
  NAND2xp33_ASAP7_75t_R  g0125( .A (x11), .B (x139), .Y (n607) );
  NOR2xp33_ASAP7_75t_R   g0126( .A (x12), .B (x140), .Y (n613) );
  NAND2xp33_ASAP7_75t_R  g0127( .A (n269), .B (n397), .Y (n605) );
  OAI21xp33_ASAP7_75t_R  g0128( .A1 (n597), .A2 (n601), .B (n605), .Y (n611) );
  AOI21xp33_ASAP7_75t_R  g0129( .A1 (n607), .B (n613), .A2 (n611), .Y (n619) );
  NOR2xp33_ASAP7_75t_R   g0130( .A (n615), .B (n619), .Y (n621) );
  INVx1_ASAP7_75t_R      g0131( .A (x13), .Y (n271) );
  XNOR2xp5_ASAP7_75t_R   g0132( .A (n271), .B (x141), .Y (n626) );
  XNOR2xp5_ASAP7_75t_R   g0133( .A (n621), .B (n626), .Y (y13) );
  INVx1_ASAP7_75t_R      g0134( .A (x141), .Y (n399) );
  NOR2xp33_ASAP7_75t_R   g0135( .A (n271), .B (n399), .Y (n624) );
  NAND2xp33_ASAP7_75t_R  g0136( .A (x12), .B (x140), .Y (n616) );
  NOR2xp33_ASAP7_75t_R   g0137( .A (x13), .B (x141), .Y (n622) );
  NAND2xp33_ASAP7_75t_R  g0138( .A (n270), .B (n398), .Y (n614) );
  OAI21xp33_ASAP7_75t_R  g0139( .A1 (n606), .A2 (n610), .B (n614), .Y (n620) );
  AOI21xp33_ASAP7_75t_R  g0140( .A1 (n616), .B (n622), .A2 (n620), .Y (n628) );
  NOR2xp33_ASAP7_75t_R   g0141( .A (n624), .B (n628), .Y (n630) );
  INVx1_ASAP7_75t_R      g0142( .A (x14), .Y (n272) );
  XNOR2xp5_ASAP7_75t_R   g0143( .A (n272), .B (x142), .Y (n635) );
  XNOR2xp5_ASAP7_75t_R   g0144( .A (n630), .B (n635), .Y (y14) );
  INVx1_ASAP7_75t_R      g0145( .A (x142), .Y (n400) );
  NOR2xp33_ASAP7_75t_R   g0146( .A (n272), .B (n400), .Y (n633) );
  NAND2xp33_ASAP7_75t_R  g0147( .A (x13), .B (x141), .Y (n625) );
  NOR2xp33_ASAP7_75t_R   g0148( .A (x14), .B (x142), .Y (n631) );
  NAND2xp33_ASAP7_75t_R  g0149( .A (n271), .B (n399), .Y (n623) );
  OAI21xp33_ASAP7_75t_R  g0150( .A1 (n615), .A2 (n619), .B (n623), .Y (n629) );
  AOI21xp33_ASAP7_75t_R  g0151( .A1 (n625), .B (n631), .A2 (n629), .Y (n637) );
  NOR2xp33_ASAP7_75t_R   g0152( .A (n633), .B (n637), .Y (n639) );
  INVx1_ASAP7_75t_R      g0153( .A (x15), .Y (n273) );
  XNOR2xp5_ASAP7_75t_R   g0154( .A (n273), .B (x143), .Y (n644) );
  XNOR2xp5_ASAP7_75t_R   g0155( .A (n639), .B (n644), .Y (y15) );
  INVx1_ASAP7_75t_R      g0156( .A (x143), .Y (n401) );
  NOR2xp33_ASAP7_75t_R   g0157( .A (n273), .B (n401), .Y (n642) );
  NAND2xp33_ASAP7_75t_R  g0158( .A (x14), .B (x142), .Y (n634) );
  NOR2xp33_ASAP7_75t_R   g0159( .A (x15), .B (x143), .Y (n640) );
  NAND2xp33_ASAP7_75t_R  g0160( .A (n272), .B (n400), .Y (n632) );
  OAI21xp33_ASAP7_75t_R  g0161( .A1 (n624), .A2 (n628), .B (n632), .Y (n638) );
  AOI21xp33_ASAP7_75t_R  g0162( .A1 (n634), .B (n640), .A2 (n638), .Y (n646) );
  NOR2xp33_ASAP7_75t_R   g0163( .A (n642), .B (n646), .Y (n648) );
  INVx1_ASAP7_75t_R      g0164( .A (x16), .Y (n274) );
  XNOR2xp5_ASAP7_75t_R   g0165( .A (n274), .B (x144), .Y (n653) );
  XNOR2xp5_ASAP7_75t_R   g0166( .A (n648), .B (n653), .Y (y16) );
  INVx1_ASAP7_75t_R      g0167( .A (x144), .Y (n402) );
  NOR2xp33_ASAP7_75t_R   g0168( .A (n274), .B (n402), .Y (n651) );
  NAND2xp33_ASAP7_75t_R  g0169( .A (x15), .B (x143), .Y (n643) );
  NOR2xp33_ASAP7_75t_R   g0170( .A (x16), .B (x144), .Y (n649) );
  NAND2xp33_ASAP7_75t_R  g0171( .A (n273), .B (n401), .Y (n641) );
  OAI21xp33_ASAP7_75t_R  g0172( .A1 (n633), .A2 (n637), .B (n641), .Y (n647) );
  AOI21xp33_ASAP7_75t_R  g0173( .A1 (n643), .B (n649), .A2 (n647), .Y (n655) );
  NOR2xp33_ASAP7_75t_R   g0174( .A (n651), .B (n655), .Y (n657) );
  INVx1_ASAP7_75t_R      g0175( .A (x17), .Y (n275) );
  XNOR2xp5_ASAP7_75t_R   g0176( .A (n275), .B (x145), .Y (n662) );
  XNOR2xp5_ASAP7_75t_R   g0177( .A (n657), .B (n662), .Y (y17) );
  INVx1_ASAP7_75t_R      g0178( .A (x145), .Y (n403) );
  NOR2xp33_ASAP7_75t_R   g0179( .A (n275), .B (n403), .Y (n660) );
  NAND2xp33_ASAP7_75t_R  g0180( .A (x16), .B (x144), .Y (n652) );
  NOR2xp33_ASAP7_75t_R   g0181( .A (x17), .B (x145), .Y (n658) );
  NAND2xp33_ASAP7_75t_R  g0182( .A (n274), .B (n402), .Y (n650) );
  OAI21xp33_ASAP7_75t_R  g0183( .A1 (n642), .A2 (n646), .B (n650), .Y (n656) );
  AOI21xp33_ASAP7_75t_R  g0184( .A1 (n652), .B (n658), .A2 (n656), .Y (n664) );
  NOR2xp33_ASAP7_75t_R   g0185( .A (n660), .B (n664), .Y (n666) );
  INVx1_ASAP7_75t_R      g0186( .A (x18), .Y (n276) );
  XNOR2xp5_ASAP7_75t_R   g0187( .A (n276), .B (x146), .Y (n671) );
  XNOR2xp5_ASAP7_75t_R   g0188( .A (n666), .B (n671), .Y (y18) );
  INVx1_ASAP7_75t_R      g0189( .A (x146), .Y (n404) );
  NOR2xp33_ASAP7_75t_R   g0190( .A (n276), .B (n404), .Y (n669) );
  NAND2xp33_ASAP7_75t_R  g0191( .A (x17), .B (x145), .Y (n661) );
  NOR2xp33_ASAP7_75t_R   g0192( .A (x18), .B (x146), .Y (n667) );
  NAND2xp33_ASAP7_75t_R  g0193( .A (n275), .B (n403), .Y (n659) );
  OAI21xp33_ASAP7_75t_R  g0194( .A1 (n651), .A2 (n655), .B (n659), .Y (n665) );
  AOI21xp33_ASAP7_75t_R  g0195( .A1 (n661), .B (n667), .A2 (n665), .Y (n673) );
  NOR2xp33_ASAP7_75t_R   g0196( .A (n669), .B (n673), .Y (n675) );
  INVx1_ASAP7_75t_R      g0197( .A (x19), .Y (n277) );
  XNOR2xp5_ASAP7_75t_R   g0198( .A (n277), .B (x147), .Y (n680) );
  XNOR2xp5_ASAP7_75t_R   g0199( .A (n675), .B (n680), .Y (y19) );
  INVx1_ASAP7_75t_R      g0200( .A (x147), .Y (n405) );
  NOR2xp33_ASAP7_75t_R   g0201( .A (n277), .B (n405), .Y (n678) );
  NAND2xp33_ASAP7_75t_R  g0202( .A (x18), .B (x146), .Y (n670) );
  NOR2xp33_ASAP7_75t_R   g0203( .A (x19), .B (x147), .Y (n676) );
  NAND2xp33_ASAP7_75t_R  g0204( .A (n276), .B (n404), .Y (n668) );
  OAI21xp33_ASAP7_75t_R  g0205( .A1 (n660), .A2 (n664), .B (n668), .Y (n674) );
  AOI21xp33_ASAP7_75t_R  g0206( .A1 (n670), .B (n676), .A2 (n674), .Y (n682) );
  NOR2xp33_ASAP7_75t_R   g0207( .A (n678), .B (n682), .Y (n684) );
  INVx1_ASAP7_75t_R      g0208( .A (x20), .Y (n278) );
  XNOR2xp5_ASAP7_75t_R   g0209( .A (n278), .B (x148), .Y (n689) );
  XNOR2xp5_ASAP7_75t_R   g0210( .A (n684), .B (n689), .Y (y20) );
  INVx1_ASAP7_75t_R      g0211( .A (x148), .Y (n406) );
  NOR2xp33_ASAP7_75t_R   g0212( .A (n278), .B (n406), .Y (n687) );
  NAND2xp33_ASAP7_75t_R  g0213( .A (x19), .B (x147), .Y (n679) );
  NOR2xp33_ASAP7_75t_R   g0214( .A (x20), .B (x148), .Y (n685) );
  NAND2xp33_ASAP7_75t_R  g0215( .A (n277), .B (n405), .Y (n677) );
  OAI21xp33_ASAP7_75t_R  g0216( .A1 (n669), .A2 (n673), .B (n677), .Y (n683) );
  AOI21xp33_ASAP7_75t_R  g0217( .A1 (n679), .B (n685), .A2 (n683), .Y (n691) );
  NOR2xp33_ASAP7_75t_R   g0218( .A (n687), .B (n691), .Y (n693) );
  INVx1_ASAP7_75t_R      g0219( .A (x21), .Y (n279) );
  XNOR2xp5_ASAP7_75t_R   g0220( .A (n279), .B (x149), .Y (n698) );
  XNOR2xp5_ASAP7_75t_R   g0221( .A (n693), .B (n698), .Y (y21) );
  INVx1_ASAP7_75t_R      g0222( .A (x149), .Y (n407) );
  NOR2xp33_ASAP7_75t_R   g0223( .A (n279), .B (n407), .Y (n696) );
  NAND2xp33_ASAP7_75t_R  g0224( .A (x20), .B (x148), .Y (n688) );
  NOR2xp33_ASAP7_75t_R   g0225( .A (x21), .B (x149), .Y (n694) );
  NAND2xp33_ASAP7_75t_R  g0226( .A (n278), .B (n406), .Y (n686) );
  OAI21xp33_ASAP7_75t_R  g0227( .A1 (n678), .A2 (n682), .B (n686), .Y (n692) );
  AOI21xp33_ASAP7_75t_R  g0228( .A1 (n688), .B (n694), .A2 (n692), .Y (n700) );
  NOR2xp33_ASAP7_75t_R   g0229( .A (n696), .B (n700), .Y (n702) );
  INVx1_ASAP7_75t_R      g0230( .A (x22), .Y (n280) );
  XNOR2xp5_ASAP7_75t_R   g0231( .A (n280), .B (x150), .Y (n707) );
  XNOR2xp5_ASAP7_75t_R   g0232( .A (n702), .B (n707), .Y (y22) );
  INVx1_ASAP7_75t_R      g0233( .A (x150), .Y (n408) );
  NOR2xp33_ASAP7_75t_R   g0234( .A (n280), .B (n408), .Y (n705) );
  NAND2xp33_ASAP7_75t_R  g0235( .A (x21), .B (x149), .Y (n697) );
  NOR2xp33_ASAP7_75t_R   g0236( .A (x22), .B (x150), .Y (n703) );
  NAND2xp33_ASAP7_75t_R  g0237( .A (n279), .B (n407), .Y (n695) );
  OAI21xp33_ASAP7_75t_R  g0238( .A1 (n687), .A2 (n691), .B (n695), .Y (n701) );
  AOI21xp33_ASAP7_75t_R  g0239( .A1 (n697), .B (n703), .A2 (n701), .Y (n709) );
  NOR2xp33_ASAP7_75t_R   g0240( .A (n705), .B (n709), .Y (n711) );
  INVx1_ASAP7_75t_R      g0241( .A (x23), .Y (n281) );
  XNOR2xp5_ASAP7_75t_R   g0242( .A (n281), .B (x151), .Y (n716) );
  XNOR2xp5_ASAP7_75t_R   g0243( .A (n711), .B (n716), .Y (y23) );
  INVx1_ASAP7_75t_R      g0244( .A (x151), .Y (n409) );
  NOR2xp33_ASAP7_75t_R   g0245( .A (n281), .B (n409), .Y (n714) );
  NAND2xp33_ASAP7_75t_R  g0246( .A (x22), .B (x150), .Y (n706) );
  NOR2xp33_ASAP7_75t_R   g0247( .A (x23), .B (x151), .Y (n712) );
  NAND2xp33_ASAP7_75t_R  g0248( .A (n280), .B (n408), .Y (n704) );
  OAI21xp33_ASAP7_75t_R  g0249( .A1 (n696), .A2 (n700), .B (n704), .Y (n710) );
  AOI21xp33_ASAP7_75t_R  g0250( .A1 (n706), .B (n712), .A2 (n710), .Y (n718) );
  NOR2xp33_ASAP7_75t_R   g0251( .A (n714), .B (n718), .Y (n720) );
  INVx1_ASAP7_75t_R      g0252( .A (x24), .Y (n282) );
  XNOR2xp5_ASAP7_75t_R   g0253( .A (n282), .B (x152), .Y (n725) );
  XNOR2xp5_ASAP7_75t_R   g0254( .A (n720), .B (n725), .Y (y24) );
  INVx1_ASAP7_75t_R      g0255( .A (x152), .Y (n410) );
  NOR2xp33_ASAP7_75t_R   g0256( .A (n282), .B (n410), .Y (n723) );
  NAND2xp33_ASAP7_75t_R  g0257( .A (x23), .B (x151), .Y (n715) );
  NOR2xp33_ASAP7_75t_R   g0258( .A (x24), .B (x152), .Y (n721) );
  NAND2xp33_ASAP7_75t_R  g0259( .A (n281), .B (n409), .Y (n713) );
  OAI21xp33_ASAP7_75t_R  g0260( .A1 (n705), .A2 (n709), .B (n713), .Y (n719) );
  AOI21xp33_ASAP7_75t_R  g0261( .A1 (n715), .B (n721), .A2 (n719), .Y (n727) );
  NOR2xp33_ASAP7_75t_R   g0262( .A (n723), .B (n727), .Y (n729) );
  INVx1_ASAP7_75t_R      g0263( .A (x25), .Y (n283) );
  XNOR2xp5_ASAP7_75t_R   g0264( .A (n283), .B (x153), .Y (n734) );
  XNOR2xp5_ASAP7_75t_R   g0265( .A (n729), .B (n734), .Y (y25) );
  INVx1_ASAP7_75t_R      g0266( .A (x153), .Y (n411) );
  NOR2xp33_ASAP7_75t_R   g0267( .A (n283), .B (n411), .Y (n732) );
  NAND2xp33_ASAP7_75t_R  g0268( .A (x24), .B (x152), .Y (n724) );
  NOR2xp33_ASAP7_75t_R   g0269( .A (x25), .B (x153), .Y (n730) );
  NAND2xp33_ASAP7_75t_R  g0270( .A (n282), .B (n410), .Y (n722) );
  OAI21xp33_ASAP7_75t_R  g0271( .A1 (n714), .A2 (n718), .B (n722), .Y (n728) );
  AOI21xp33_ASAP7_75t_R  g0272( .A1 (n724), .B (n730), .A2 (n728), .Y (n736) );
  NOR2xp33_ASAP7_75t_R   g0273( .A (n732), .B (n736), .Y (n738) );
  INVx1_ASAP7_75t_R      g0274( .A (x26), .Y (n284) );
  XNOR2xp5_ASAP7_75t_R   g0275( .A (n284), .B (x154), .Y (n743) );
  XNOR2xp5_ASAP7_75t_R   g0276( .A (n738), .B (n743), .Y (y26) );
  INVx1_ASAP7_75t_R      g0277( .A (x154), .Y (n412) );
  NOR2xp33_ASAP7_75t_R   g0278( .A (n284), .B (n412), .Y (n741) );
  NAND2xp33_ASAP7_75t_R  g0279( .A (x25), .B (x153), .Y (n733) );
  NOR2xp33_ASAP7_75t_R   g0280( .A (x26), .B (x154), .Y (n739) );
  NAND2xp33_ASAP7_75t_R  g0281( .A (n283), .B (n411), .Y (n731) );
  OAI21xp33_ASAP7_75t_R  g0282( .A1 (n723), .A2 (n727), .B (n731), .Y (n737) );
  AOI21xp33_ASAP7_75t_R  g0283( .A1 (n733), .B (n739), .A2 (n737), .Y (n745) );
  NOR2xp33_ASAP7_75t_R   g0284( .A (n741), .B (n745), .Y (n747) );
  INVx1_ASAP7_75t_R      g0285( .A (x27), .Y (n285) );
  XNOR2xp5_ASAP7_75t_R   g0286( .A (n285), .B (x155), .Y (n752) );
  XNOR2xp5_ASAP7_75t_R   g0287( .A (n747), .B (n752), .Y (y27) );
  INVx1_ASAP7_75t_R      g0288( .A (x155), .Y (n413) );
  NOR2xp33_ASAP7_75t_R   g0289( .A (n285), .B (n413), .Y (n750) );
  NAND2xp33_ASAP7_75t_R  g0290( .A (x26), .B (x154), .Y (n742) );
  NOR2xp33_ASAP7_75t_R   g0291( .A (x27), .B (x155), .Y (n748) );
  NAND2xp33_ASAP7_75t_R  g0292( .A (n284), .B (n412), .Y (n740) );
  OAI21xp33_ASAP7_75t_R  g0293( .A1 (n732), .A2 (n736), .B (n740), .Y (n746) );
  AOI21xp33_ASAP7_75t_R  g0294( .A1 (n742), .B (n748), .A2 (n746), .Y (n754) );
  NOR2xp33_ASAP7_75t_R   g0295( .A (n750), .B (n754), .Y (n756) );
  INVx1_ASAP7_75t_R      g0296( .A (x28), .Y (n286) );
  XNOR2xp5_ASAP7_75t_R   g0297( .A (n286), .B (x156), .Y (n761) );
  XNOR2xp5_ASAP7_75t_R   g0298( .A (n756), .B (n761), .Y (y28) );
  INVx1_ASAP7_75t_R      g0299( .A (x156), .Y (n414) );
  NOR2xp33_ASAP7_75t_R   g0300( .A (n286), .B (n414), .Y (n759) );
  NAND2xp33_ASAP7_75t_R  g0301( .A (x27), .B (x155), .Y (n751) );
  NOR2xp33_ASAP7_75t_R   g0302( .A (x28), .B (x156), .Y (n757) );
  NAND2xp33_ASAP7_75t_R  g0303( .A (n285), .B (n413), .Y (n749) );
  OAI21xp33_ASAP7_75t_R  g0304( .A1 (n741), .A2 (n745), .B (n749), .Y (n755) );
  AOI21xp33_ASAP7_75t_R  g0305( .A1 (n751), .B (n757), .A2 (n755), .Y (n763) );
  NOR2xp33_ASAP7_75t_R   g0306( .A (n759), .B (n763), .Y (n765) );
  INVx1_ASAP7_75t_R      g0307( .A (x29), .Y (n287) );
  XNOR2xp5_ASAP7_75t_R   g0308( .A (n287), .B (x157), .Y (n770) );
  XNOR2xp5_ASAP7_75t_R   g0309( .A (n765), .B (n770), .Y (y29) );
  INVx1_ASAP7_75t_R      g0310( .A (x157), .Y (n415) );
  NOR2xp33_ASAP7_75t_R   g0311( .A (n287), .B (n415), .Y (n768) );
  NAND2xp33_ASAP7_75t_R  g0312( .A (x28), .B (x156), .Y (n760) );
  NOR2xp33_ASAP7_75t_R   g0313( .A (x29), .B (x157), .Y (n766) );
  NAND2xp33_ASAP7_75t_R  g0314( .A (n286), .B (n414), .Y (n758) );
  OAI21xp33_ASAP7_75t_R  g0315( .A1 (n750), .A2 (n754), .B (n758), .Y (n764) );
  AOI21xp33_ASAP7_75t_R  g0316( .A1 (n760), .B (n766), .A2 (n764), .Y (n772) );
  NOR2xp33_ASAP7_75t_R   g0317( .A (n768), .B (n772), .Y (n774) );
  INVx1_ASAP7_75t_R      g0318( .A (x30), .Y (n288) );
  XNOR2xp5_ASAP7_75t_R   g0319( .A (n288), .B (x158), .Y (n779) );
  XNOR2xp5_ASAP7_75t_R   g0320( .A (n774), .B (n779), .Y (y30) );
  INVx1_ASAP7_75t_R      g0321( .A (x158), .Y (n416) );
  NOR2xp33_ASAP7_75t_R   g0322( .A (n288), .B (n416), .Y (n777) );
  NAND2xp33_ASAP7_75t_R  g0323( .A (x29), .B (x157), .Y (n769) );
  NOR2xp33_ASAP7_75t_R   g0324( .A (x30), .B (x158), .Y (n775) );
  NAND2xp33_ASAP7_75t_R  g0325( .A (n287), .B (n415), .Y (n767) );
  OAI21xp33_ASAP7_75t_R  g0326( .A1 (n759), .A2 (n763), .B (n767), .Y (n773) );
  AOI21xp33_ASAP7_75t_R  g0327( .A1 (n769), .B (n775), .A2 (n773), .Y (n781) );
  NOR2xp33_ASAP7_75t_R   g0328( .A (n777), .B (n781), .Y (n783) );
  INVx1_ASAP7_75t_R      g0329( .A (x31), .Y (n289) );
  XNOR2xp5_ASAP7_75t_R   g0330( .A (n289), .B (x159), .Y (n788) );
  XNOR2xp5_ASAP7_75t_R   g0331( .A (n783), .B (n788), .Y (y31) );
  INVx1_ASAP7_75t_R      g0332( .A (x159), .Y (n417) );
  NOR2xp33_ASAP7_75t_R   g0333( .A (n289), .B (n417), .Y (n786) );
  NAND2xp33_ASAP7_75t_R  g0334( .A (x30), .B (x158), .Y (n778) );
  NOR2xp33_ASAP7_75t_R   g0335( .A (x31), .B (x159), .Y (n784) );
  NAND2xp33_ASAP7_75t_R  g0336( .A (n288), .B (n416), .Y (n776) );
  OAI21xp33_ASAP7_75t_R  g0337( .A1 (n768), .A2 (n772), .B (n776), .Y (n782) );
  AOI21xp33_ASAP7_75t_R  g0338( .A1 (n778), .B (n784), .A2 (n782), .Y (n790) );
  NOR2xp33_ASAP7_75t_R   g0339( .A (n786), .B (n790), .Y (n792) );
  INVx1_ASAP7_75t_R      g0340( .A (x32), .Y (n290) );
  XNOR2xp5_ASAP7_75t_R   g0341( .A (n290), .B (x160), .Y (n797) );
  XNOR2xp5_ASAP7_75t_R   g0342( .A (n792), .B (n797), .Y (y32) );
  INVx1_ASAP7_75t_R      g0343( .A (x160), .Y (n418) );
  NOR2xp33_ASAP7_75t_R   g0344( .A (n290), .B (n418), .Y (n795) );
  NAND2xp33_ASAP7_75t_R  g0345( .A (x31), .B (x159), .Y (n787) );
  NOR2xp33_ASAP7_75t_R   g0346( .A (x32), .B (x160), .Y (n793) );
  NAND2xp33_ASAP7_75t_R  g0347( .A (n289), .B (n417), .Y (n785) );
  OAI21xp33_ASAP7_75t_R  g0348( .A1 (n777), .A2 (n781), .B (n785), .Y (n791) );
  AOI21xp33_ASAP7_75t_R  g0349( .A1 (n787), .B (n793), .A2 (n791), .Y (n799) );
  NOR2xp33_ASAP7_75t_R   g0350( .A (n795), .B (n799), .Y (n801) );
  INVx1_ASAP7_75t_R      g0351( .A (x33), .Y (n291) );
  XNOR2xp5_ASAP7_75t_R   g0352( .A (n291), .B (x161), .Y (n806) );
  XNOR2xp5_ASAP7_75t_R   g0353( .A (n801), .B (n806), .Y (y33) );
  INVx1_ASAP7_75t_R      g0354( .A (x161), .Y (n419) );
  NOR2xp33_ASAP7_75t_R   g0355( .A (n291), .B (n419), .Y (n804) );
  NAND2xp33_ASAP7_75t_R  g0356( .A (x32), .B (x160), .Y (n796) );
  NOR2xp33_ASAP7_75t_R   g0357( .A (x33), .B (x161), .Y (n802) );
  NAND2xp33_ASAP7_75t_R  g0358( .A (n290), .B (n418), .Y (n794) );
  OAI21xp33_ASAP7_75t_R  g0359( .A1 (n786), .A2 (n790), .B (n794), .Y (n800) );
  AOI21xp33_ASAP7_75t_R  g0360( .A1 (n796), .B (n802), .A2 (n800), .Y (n808) );
  NOR2xp33_ASAP7_75t_R   g0361( .A (n804), .B (n808), .Y (n810) );
  INVx1_ASAP7_75t_R      g0362( .A (x34), .Y (n292) );
  XNOR2xp5_ASAP7_75t_R   g0363( .A (n292), .B (x162), .Y (n815) );
  XNOR2xp5_ASAP7_75t_R   g0364( .A (n810), .B (n815), .Y (y34) );
  INVx1_ASAP7_75t_R      g0365( .A (x162), .Y (n420) );
  NOR2xp33_ASAP7_75t_R   g0366( .A (n292), .B (n420), .Y (n813) );
  NAND2xp33_ASAP7_75t_R  g0367( .A (x33), .B (x161), .Y (n805) );
  NOR2xp33_ASAP7_75t_R   g0368( .A (x34), .B (x162), .Y (n811) );
  NAND2xp33_ASAP7_75t_R  g0369( .A (n291), .B (n419), .Y (n803) );
  OAI21xp33_ASAP7_75t_R  g0370( .A1 (n795), .A2 (n799), .B (n803), .Y (n809) );
  AOI21xp33_ASAP7_75t_R  g0371( .A1 (n805), .B (n811), .A2 (n809), .Y (n817) );
  NOR2xp33_ASAP7_75t_R   g0372( .A (n813), .B (n817), .Y (n819) );
  INVx1_ASAP7_75t_R      g0373( .A (x35), .Y (n293) );
  XNOR2xp5_ASAP7_75t_R   g0374( .A (n293), .B (x163), .Y (n824) );
  XNOR2xp5_ASAP7_75t_R   g0375( .A (n819), .B (n824), .Y (y35) );
  INVx1_ASAP7_75t_R      g0376( .A (x163), .Y (n421) );
  NOR2xp33_ASAP7_75t_R   g0377( .A (n293), .B (n421), .Y (n822) );
  NAND2xp33_ASAP7_75t_R  g0378( .A (x34), .B (x162), .Y (n814) );
  NOR2xp33_ASAP7_75t_R   g0379( .A (x35), .B (x163), .Y (n820) );
  NAND2xp33_ASAP7_75t_R  g0380( .A (n292), .B (n420), .Y (n812) );
  OAI21xp33_ASAP7_75t_R  g0381( .A1 (n804), .A2 (n808), .B (n812), .Y (n818) );
  AOI21xp33_ASAP7_75t_R  g0382( .A1 (n814), .B (n820), .A2 (n818), .Y (n826) );
  NOR2xp33_ASAP7_75t_R   g0383( .A (n822), .B (n826), .Y (n828) );
  INVx1_ASAP7_75t_R      g0384( .A (x36), .Y (n294) );
  XNOR2xp5_ASAP7_75t_R   g0385( .A (n294), .B (x164), .Y (n833) );
  XNOR2xp5_ASAP7_75t_R   g0386( .A (n828), .B (n833), .Y (y36) );
  INVx1_ASAP7_75t_R      g0387( .A (x164), .Y (n422) );
  NOR2xp33_ASAP7_75t_R   g0388( .A (n294), .B (n422), .Y (n831) );
  NAND2xp33_ASAP7_75t_R  g0389( .A (x35), .B (x163), .Y (n823) );
  NOR2xp33_ASAP7_75t_R   g0390( .A (x36), .B (x164), .Y (n829) );
  NAND2xp33_ASAP7_75t_R  g0391( .A (n293), .B (n421), .Y (n821) );
  OAI21xp33_ASAP7_75t_R  g0392( .A1 (n813), .A2 (n817), .B (n821), .Y (n827) );
  AOI21xp33_ASAP7_75t_R  g0393( .A1 (n823), .B (n829), .A2 (n827), .Y (n835) );
  NOR2xp33_ASAP7_75t_R   g0394( .A (n831), .B (n835), .Y (n837) );
  INVx1_ASAP7_75t_R      g0395( .A (x37), .Y (n295) );
  XNOR2xp5_ASAP7_75t_R   g0396( .A (n295), .B (x165), .Y (n842) );
  XNOR2xp5_ASAP7_75t_R   g0397( .A (n837), .B (n842), .Y (y37) );
  INVx1_ASAP7_75t_R      g0398( .A (x165), .Y (n423) );
  NOR2xp33_ASAP7_75t_R   g0399( .A (n295), .B (n423), .Y (n840) );
  NAND2xp33_ASAP7_75t_R  g0400( .A (x36), .B (x164), .Y (n832) );
  NOR2xp33_ASAP7_75t_R   g0401( .A (x37), .B (x165), .Y (n838) );
  NAND2xp33_ASAP7_75t_R  g0402( .A (n294), .B (n422), .Y (n830) );
  OAI21xp33_ASAP7_75t_R  g0403( .A1 (n822), .A2 (n826), .B (n830), .Y (n836) );
  AOI21xp33_ASAP7_75t_R  g0404( .A1 (n832), .B (n838), .A2 (n836), .Y (n844) );
  NOR2xp33_ASAP7_75t_R   g0405( .A (n840), .B (n844), .Y (n846) );
  INVx1_ASAP7_75t_R      g0406( .A (x38), .Y (n296) );
  XNOR2xp5_ASAP7_75t_R   g0407( .A (n296), .B (x166), .Y (n851) );
  XNOR2xp5_ASAP7_75t_R   g0408( .A (n846), .B (n851), .Y (y38) );
  INVx1_ASAP7_75t_R      g0409( .A (x166), .Y (n424) );
  NOR2xp33_ASAP7_75t_R   g0410( .A (n296), .B (n424), .Y (n849) );
  NAND2xp33_ASAP7_75t_R  g0411( .A (x37), .B (x165), .Y (n841) );
  NOR2xp33_ASAP7_75t_R   g0412( .A (x38), .B (x166), .Y (n847) );
  NAND2xp33_ASAP7_75t_R  g0413( .A (n295), .B (n423), .Y (n839) );
  OAI21xp33_ASAP7_75t_R  g0414( .A1 (n831), .A2 (n835), .B (n839), .Y (n845) );
  AOI21xp33_ASAP7_75t_R  g0415( .A1 (n841), .B (n847), .A2 (n845), .Y (n853) );
  NOR2xp33_ASAP7_75t_R   g0416( .A (n849), .B (n853), .Y (n855) );
  INVx1_ASAP7_75t_R      g0417( .A (x39), .Y (n297) );
  XNOR2xp5_ASAP7_75t_R   g0418( .A (n297), .B (x167), .Y (n860) );
  XNOR2xp5_ASAP7_75t_R   g0419( .A (n855), .B (n860), .Y (y39) );
  INVx1_ASAP7_75t_R      g0420( .A (x167), .Y (n425) );
  NOR2xp33_ASAP7_75t_R   g0421( .A (n297), .B (n425), .Y (n858) );
  NAND2xp33_ASAP7_75t_R  g0422( .A (x38), .B (x166), .Y (n850) );
  NOR2xp33_ASAP7_75t_R   g0423( .A (x39), .B (x167), .Y (n856) );
  NAND2xp33_ASAP7_75t_R  g0424( .A (n296), .B (n424), .Y (n848) );
  OAI21xp33_ASAP7_75t_R  g0425( .A1 (n840), .A2 (n844), .B (n848), .Y (n854) );
  AOI21xp33_ASAP7_75t_R  g0426( .A1 (n850), .B (n856), .A2 (n854), .Y (n862) );
  NOR2xp33_ASAP7_75t_R   g0427( .A (n858), .B (n862), .Y (n864) );
  INVx1_ASAP7_75t_R      g0428( .A (x40), .Y (n298) );
  XNOR2xp5_ASAP7_75t_R   g0429( .A (n298), .B (x168), .Y (n869) );
  XNOR2xp5_ASAP7_75t_R   g0430( .A (n864), .B (n869), .Y (y40) );
  INVx1_ASAP7_75t_R      g0431( .A (x168), .Y (n426) );
  NOR2xp33_ASAP7_75t_R   g0432( .A (n298), .B (n426), .Y (n867) );
  NAND2xp33_ASAP7_75t_R  g0433( .A (x39), .B (x167), .Y (n859) );
  NOR2xp33_ASAP7_75t_R   g0434( .A (x40), .B (x168), .Y (n865) );
  NAND2xp33_ASAP7_75t_R  g0435( .A (n297), .B (n425), .Y (n857) );
  OAI21xp33_ASAP7_75t_R  g0436( .A1 (n849), .A2 (n853), .B (n857), .Y (n863) );
  AOI21xp33_ASAP7_75t_R  g0437( .A1 (n859), .B (n865), .A2 (n863), .Y (n871) );
  NOR2xp33_ASAP7_75t_R   g0438( .A (n867), .B (n871), .Y (n873) );
  INVx1_ASAP7_75t_R      g0439( .A (x41), .Y (n299) );
  XNOR2xp5_ASAP7_75t_R   g0440( .A (n299), .B (x169), .Y (n878) );
  XNOR2xp5_ASAP7_75t_R   g0441( .A (n873), .B (n878), .Y (y41) );
  INVx1_ASAP7_75t_R      g0442( .A (x169), .Y (n427) );
  NOR2xp33_ASAP7_75t_R   g0443( .A (n299), .B (n427), .Y (n876) );
  NAND2xp33_ASAP7_75t_R  g0444( .A (x40), .B (x168), .Y (n868) );
  NOR2xp33_ASAP7_75t_R   g0445( .A (x41), .B (x169), .Y (n874) );
  NAND2xp33_ASAP7_75t_R  g0446( .A (n298), .B (n426), .Y (n866) );
  OAI21xp33_ASAP7_75t_R  g0447( .A1 (n858), .A2 (n862), .B (n866), .Y (n872) );
  AOI21xp33_ASAP7_75t_R  g0448( .A1 (n868), .B (n874), .A2 (n872), .Y (n880) );
  NOR2xp33_ASAP7_75t_R   g0449( .A (n876), .B (n880), .Y (n882) );
  INVx1_ASAP7_75t_R      g0450( .A (x42), .Y (n300) );
  XNOR2xp5_ASAP7_75t_R   g0451( .A (n300), .B (x170), .Y (n887) );
  XNOR2xp5_ASAP7_75t_R   g0452( .A (n882), .B (n887), .Y (y42) );
  INVx1_ASAP7_75t_R      g0453( .A (x170), .Y (n428) );
  NOR2xp33_ASAP7_75t_R   g0454( .A (n300), .B (n428), .Y (n885) );
  NAND2xp33_ASAP7_75t_R  g0455( .A (x41), .B (x169), .Y (n877) );
  NOR2xp33_ASAP7_75t_R   g0456( .A (x42), .B (x170), .Y (n883) );
  NAND2xp33_ASAP7_75t_R  g0457( .A (n299), .B (n427), .Y (n875) );
  OAI21xp33_ASAP7_75t_R  g0458( .A1 (n867), .A2 (n871), .B (n875), .Y (n881) );
  AOI21xp33_ASAP7_75t_R  g0459( .A1 (n877), .B (n883), .A2 (n881), .Y (n889) );
  NOR2xp33_ASAP7_75t_R   g0460( .A (n885), .B (n889), .Y (n891) );
  INVx1_ASAP7_75t_R      g0461( .A (x43), .Y (n301) );
  XNOR2xp5_ASAP7_75t_R   g0462( .A (n301), .B (x171), .Y (n896) );
  XNOR2xp5_ASAP7_75t_R   g0463( .A (n891), .B (n896), .Y (y43) );
  INVx1_ASAP7_75t_R      g0464( .A (x171), .Y (n429) );
  NOR2xp33_ASAP7_75t_R   g0465( .A (n301), .B (n429), .Y (n894) );
  NAND2xp33_ASAP7_75t_R  g0466( .A (x42), .B (x170), .Y (n886) );
  NOR2xp33_ASAP7_75t_R   g0467( .A (x43), .B (x171), .Y (n892) );
  NAND2xp33_ASAP7_75t_R  g0468( .A (n300), .B (n428), .Y (n884) );
  OAI21xp33_ASAP7_75t_R  g0469( .A1 (n876), .A2 (n880), .B (n884), .Y (n890) );
  AOI21xp33_ASAP7_75t_R  g0470( .A1 (n886), .B (n892), .A2 (n890), .Y (n898) );
  NOR2xp33_ASAP7_75t_R   g0471( .A (n894), .B (n898), .Y (n900) );
  INVx1_ASAP7_75t_R      g0472( .A (x44), .Y (n302) );
  XNOR2xp5_ASAP7_75t_R   g0473( .A (n302), .B (x172), .Y (n905) );
  XNOR2xp5_ASAP7_75t_R   g0474( .A (n900), .B (n905), .Y (y44) );
  INVx1_ASAP7_75t_R      g0475( .A (x172), .Y (n430) );
  NOR2xp33_ASAP7_75t_R   g0476( .A (n302), .B (n430), .Y (n903) );
  NAND2xp33_ASAP7_75t_R  g0477( .A (x43), .B (x171), .Y (n895) );
  NOR2xp33_ASAP7_75t_R   g0478( .A (x44), .B (x172), .Y (n901) );
  NAND2xp33_ASAP7_75t_R  g0479( .A (n301), .B (n429), .Y (n893) );
  OAI21xp33_ASAP7_75t_R  g0480( .A1 (n885), .A2 (n889), .B (n893), .Y (n899) );
  AOI21xp33_ASAP7_75t_R  g0481( .A1 (n895), .B (n901), .A2 (n899), .Y (n907) );
  NOR2xp33_ASAP7_75t_R   g0482( .A (n903), .B (n907), .Y (n909) );
  INVx1_ASAP7_75t_R      g0483( .A (x45), .Y (n303) );
  XNOR2xp5_ASAP7_75t_R   g0484( .A (n303), .B (x173), .Y (n914) );
  XNOR2xp5_ASAP7_75t_R   g0485( .A (n909), .B (n914), .Y (y45) );
  INVx1_ASAP7_75t_R      g0486( .A (x173), .Y (n431) );
  NOR2xp33_ASAP7_75t_R   g0487( .A (n303), .B (n431), .Y (n912) );
  NAND2xp33_ASAP7_75t_R  g0488( .A (x44), .B (x172), .Y (n904) );
  NOR2xp33_ASAP7_75t_R   g0489( .A (x45), .B (x173), .Y (n910) );
  NAND2xp33_ASAP7_75t_R  g0490( .A (n302), .B (n430), .Y (n902) );
  OAI21xp33_ASAP7_75t_R  g0491( .A1 (n894), .A2 (n898), .B (n902), .Y (n908) );
  AOI21xp33_ASAP7_75t_R  g0492( .A1 (n904), .B (n910), .A2 (n908), .Y (n916) );
  NOR2xp33_ASAP7_75t_R   g0493( .A (n912), .B (n916), .Y (n918) );
  INVx1_ASAP7_75t_R      g0494( .A (x46), .Y (n304) );
  XNOR2xp5_ASAP7_75t_R   g0495( .A (n304), .B (x174), .Y (n923) );
  XNOR2xp5_ASAP7_75t_R   g0496( .A (n918), .B (n923), .Y (y46) );
  INVx1_ASAP7_75t_R      g0497( .A (x174), .Y (n432) );
  NOR2xp33_ASAP7_75t_R   g0498( .A (n304), .B (n432), .Y (n921) );
  NAND2xp33_ASAP7_75t_R  g0499( .A (x45), .B (x173), .Y (n913) );
  NOR2xp33_ASAP7_75t_R   g0500( .A (x46), .B (x174), .Y (n919) );
  NAND2xp33_ASAP7_75t_R  g0501( .A (n303), .B (n431), .Y (n911) );
  OAI21xp33_ASAP7_75t_R  g0502( .A1 (n903), .A2 (n907), .B (n911), .Y (n917) );
  AOI21xp33_ASAP7_75t_R  g0503( .A1 (n913), .B (n919), .A2 (n917), .Y (n925) );
  NOR2xp33_ASAP7_75t_R   g0504( .A (n921), .B (n925), .Y (n927) );
  INVx1_ASAP7_75t_R      g0505( .A (x47), .Y (n305) );
  XNOR2xp5_ASAP7_75t_R   g0506( .A (n305), .B (x175), .Y (n932) );
  XNOR2xp5_ASAP7_75t_R   g0507( .A (n927), .B (n932), .Y (y47) );
  INVx1_ASAP7_75t_R      g0508( .A (x175), .Y (n433) );
  NOR2xp33_ASAP7_75t_R   g0509( .A (n305), .B (n433), .Y (n930) );
  NAND2xp33_ASAP7_75t_R  g0510( .A (x46), .B (x174), .Y (n922) );
  NOR2xp33_ASAP7_75t_R   g0511( .A (x47), .B (x175), .Y (n928) );
  NAND2xp33_ASAP7_75t_R  g0512( .A (n304), .B (n432), .Y (n920) );
  OAI21xp33_ASAP7_75t_R  g0513( .A1 (n912), .A2 (n916), .B (n920), .Y (n926) );
  AOI21xp33_ASAP7_75t_R  g0514( .A1 (n922), .B (n928), .A2 (n926), .Y (n934) );
  NOR2xp33_ASAP7_75t_R   g0515( .A (n930), .B (n934), .Y (n936) );
  INVx1_ASAP7_75t_R      g0516( .A (x48), .Y (n306) );
  XNOR2xp5_ASAP7_75t_R   g0517( .A (n306), .B (x176), .Y (n941) );
  XNOR2xp5_ASAP7_75t_R   g0518( .A (n936), .B (n941), .Y (y48) );
  INVx1_ASAP7_75t_R      g0519( .A (x176), .Y (n434) );
  NOR2xp33_ASAP7_75t_R   g0520( .A (n306), .B (n434), .Y (n939) );
  NAND2xp33_ASAP7_75t_R  g0521( .A (x47), .B (x175), .Y (n931) );
  NOR2xp33_ASAP7_75t_R   g0522( .A (x48), .B (x176), .Y (n937) );
  NAND2xp33_ASAP7_75t_R  g0523( .A (n305), .B (n433), .Y (n929) );
  OAI21xp33_ASAP7_75t_R  g0524( .A1 (n921), .A2 (n925), .B (n929), .Y (n935) );
  AOI21xp33_ASAP7_75t_R  g0525( .A1 (n931), .B (n937), .A2 (n935), .Y (n943) );
  NOR2xp33_ASAP7_75t_R   g0526( .A (n939), .B (n943), .Y (n945) );
  INVx1_ASAP7_75t_R      g0527( .A (x49), .Y (n307) );
  XNOR2xp5_ASAP7_75t_R   g0528( .A (n307), .B (x177), .Y (n950) );
  XNOR2xp5_ASAP7_75t_R   g0529( .A (n945), .B (n950), .Y (y49) );
  INVx1_ASAP7_75t_R      g0530( .A (x177), .Y (n435) );
  NOR2xp33_ASAP7_75t_R   g0531( .A (n307), .B (n435), .Y (n948) );
  NAND2xp33_ASAP7_75t_R  g0532( .A (x48), .B (x176), .Y (n940) );
  NOR2xp33_ASAP7_75t_R   g0533( .A (x49), .B (x177), .Y (n946) );
  NAND2xp33_ASAP7_75t_R  g0534( .A (n306), .B (n434), .Y (n938) );
  OAI21xp33_ASAP7_75t_R  g0535( .A1 (n930), .A2 (n934), .B (n938), .Y (n944) );
  AOI21xp33_ASAP7_75t_R  g0536( .A1 (n940), .B (n946), .A2 (n944), .Y (n952) );
  NOR2xp33_ASAP7_75t_R   g0537( .A (n948), .B (n952), .Y (n954) );
  INVx1_ASAP7_75t_R      g0538( .A (x50), .Y (n308) );
  XNOR2xp5_ASAP7_75t_R   g0539( .A (n308), .B (x178), .Y (n959) );
  XNOR2xp5_ASAP7_75t_R   g0540( .A (n954), .B (n959), .Y (y50) );
  INVx1_ASAP7_75t_R      g0541( .A (x178), .Y (n436) );
  NOR2xp33_ASAP7_75t_R   g0542( .A (n308), .B (n436), .Y (n957) );
  NAND2xp33_ASAP7_75t_R  g0543( .A (x49), .B (x177), .Y (n949) );
  NOR2xp33_ASAP7_75t_R   g0544( .A (x50), .B (x178), .Y (n955) );
  NAND2xp33_ASAP7_75t_R  g0545( .A (n307), .B (n435), .Y (n947) );
  OAI21xp33_ASAP7_75t_R  g0546( .A1 (n939), .A2 (n943), .B (n947), .Y (n953) );
  AOI21xp33_ASAP7_75t_R  g0547( .A1 (n949), .B (n955), .A2 (n953), .Y (n961) );
  NOR2xp33_ASAP7_75t_R   g0548( .A (n957), .B (n961), .Y (n963) );
  INVx1_ASAP7_75t_R      g0549( .A (x51), .Y (n309) );
  XNOR2xp5_ASAP7_75t_R   g0550( .A (n309), .B (x179), .Y (n968) );
  XNOR2xp5_ASAP7_75t_R   g0551( .A (n963), .B (n968), .Y (y51) );
  INVx1_ASAP7_75t_R      g0552( .A (x179), .Y (n437) );
  NOR2xp33_ASAP7_75t_R   g0553( .A (n309), .B (n437), .Y (n966) );
  NAND2xp33_ASAP7_75t_R  g0554( .A (x50), .B (x178), .Y (n958) );
  NOR2xp33_ASAP7_75t_R   g0555( .A (x51), .B (x179), .Y (n964) );
  NAND2xp33_ASAP7_75t_R  g0556( .A (n308), .B (n436), .Y (n956) );
  OAI21xp33_ASAP7_75t_R  g0557( .A1 (n948), .A2 (n952), .B (n956), .Y (n962) );
  AOI21xp33_ASAP7_75t_R  g0558( .A1 (n958), .B (n964), .A2 (n962), .Y (n970) );
  NOR2xp33_ASAP7_75t_R   g0559( .A (n966), .B (n970), .Y (n972) );
  INVx1_ASAP7_75t_R      g0560( .A (x52), .Y (n310) );
  XNOR2xp5_ASAP7_75t_R   g0561( .A (n310), .B (x180), .Y (n977) );
  XNOR2xp5_ASAP7_75t_R   g0562( .A (n972), .B (n977), .Y (y52) );
  INVx1_ASAP7_75t_R      g0563( .A (x180), .Y (n438) );
  NOR2xp33_ASAP7_75t_R   g0564( .A (n310), .B (n438), .Y (n975) );
  NAND2xp33_ASAP7_75t_R  g0565( .A (x51), .B (x179), .Y (n967) );
  NOR2xp33_ASAP7_75t_R   g0566( .A (x52), .B (x180), .Y (n973) );
  NAND2xp33_ASAP7_75t_R  g0567( .A (n309), .B (n437), .Y (n965) );
  OAI21xp33_ASAP7_75t_R  g0568( .A1 (n957), .A2 (n961), .B (n965), .Y (n971) );
  AOI21xp33_ASAP7_75t_R  g0569( .A1 (n967), .B (n973), .A2 (n971), .Y (n979) );
  NOR2xp33_ASAP7_75t_R   g0570( .A (n975), .B (n979), .Y (n981) );
  INVx1_ASAP7_75t_R      g0571( .A (x53), .Y (n311) );
  XNOR2xp5_ASAP7_75t_R   g0572( .A (n311), .B (x181), .Y (n986) );
  XNOR2xp5_ASAP7_75t_R   g0573( .A (n981), .B (n986), .Y (y53) );
  INVx1_ASAP7_75t_R      g0574( .A (x181), .Y (n439) );
  NOR2xp33_ASAP7_75t_R   g0575( .A (n311), .B (n439), .Y (n984) );
  NAND2xp33_ASAP7_75t_R  g0576( .A (x52), .B (x180), .Y (n976) );
  NOR2xp33_ASAP7_75t_R   g0577( .A (x53), .B (x181), .Y (n982) );
  NAND2xp33_ASAP7_75t_R  g0578( .A (n310), .B (n438), .Y (n974) );
  OAI21xp33_ASAP7_75t_R  g0579( .A1 (n966), .A2 (n970), .B (n974), .Y (n980) );
  AOI21xp33_ASAP7_75t_R  g0580( .A1 (n976), .B (n982), .A2 (n980), .Y (n988) );
  NOR2xp33_ASAP7_75t_R   g0581( .A (n984), .B (n988), .Y (n990) );
  INVx1_ASAP7_75t_R      g0582( .A (x54), .Y (n312) );
  XNOR2xp5_ASAP7_75t_R   g0583( .A (n312), .B (x182), .Y (n995) );
  XNOR2xp5_ASAP7_75t_R   g0584( .A (n990), .B (n995), .Y (y54) );
  INVx1_ASAP7_75t_R      g0585( .A (x182), .Y (n440) );
  NOR2xp33_ASAP7_75t_R   g0586( .A (n312), .B (n440), .Y (n993) );
  NAND2xp33_ASAP7_75t_R  g0587( .A (x53), .B (x181), .Y (n985) );
  NOR2xp33_ASAP7_75t_R   g0588( .A (x54), .B (x182), .Y (n991) );
  NAND2xp33_ASAP7_75t_R  g0589( .A (n311), .B (n439), .Y (n983) );
  OAI21xp33_ASAP7_75t_R  g0590( .A1 (n975), .A2 (n979), .B (n983), .Y (n989) );
  AOI21xp33_ASAP7_75t_R  g0591( .A1 (n985), .B (n991), .A2 (n989), .Y (n997) );
  NOR2xp33_ASAP7_75t_R   g0592( .A (n993), .B (n997), .Y (n999) );
  INVx1_ASAP7_75t_R      g0593( .A (x55), .Y (n313) );
  XNOR2xp5_ASAP7_75t_R   g0594( .A (n313), .B (x183), .Y (n1004) );
  XNOR2xp5_ASAP7_75t_R   g0595( .A (n999), .B (n1004), .Y (y55) );
  INVx1_ASAP7_75t_R      g0596( .A (x183), .Y (n441) );
  NOR2xp33_ASAP7_75t_R   g0597( .A (n313), .B (n441), .Y (n1002) );
  NAND2xp33_ASAP7_75t_R  g0598( .A (x54), .B (x182), .Y (n994) );
  NOR2xp33_ASAP7_75t_R   g0599( .A (x55), .B (x183), .Y (n1000) );
  NAND2xp33_ASAP7_75t_R  g0600( .A (n312), .B (n440), .Y (n992) );
  OAI21xp33_ASAP7_75t_R  g0601( .A1 (n984), .A2 (n988), .B (n992), .Y (n998) );
  AOI21xp33_ASAP7_75t_R  g0602( .A1 (n994), .B (n1000), .A2 (n998), .Y (n1006) );
  NOR2xp33_ASAP7_75t_R   g0603( .A (n1002), .B (n1006), .Y (n1008) );
  INVx1_ASAP7_75t_R      g0604( .A (x56), .Y (n314) );
  XNOR2xp5_ASAP7_75t_R   g0605( .A (n314), .B (x184), .Y (n1013) );
  XNOR2xp5_ASAP7_75t_R   g0606( .A (n1008), .B (n1013), .Y (y56) );
  INVx1_ASAP7_75t_R      g0607( .A (x184), .Y (n442) );
  NOR2xp33_ASAP7_75t_R   g0608( .A (n314), .B (n442), .Y (n1011) );
  NAND2xp33_ASAP7_75t_R  g0609( .A (x55), .B (x183), .Y (n1003) );
  NOR2xp33_ASAP7_75t_R   g0610( .A (x56), .B (x184), .Y (n1009) );
  NAND2xp33_ASAP7_75t_R  g0611( .A (n313), .B (n441), .Y (n1001) );
  OAI21xp33_ASAP7_75t_R  g0612( .A1 (n993), .A2 (n997), .B (n1001), .Y (n1007) );
  AOI21xp33_ASAP7_75t_R  g0613( .A1 (n1003), .B (n1009), .A2 (n1007), .Y (n1015) );
  NOR2xp33_ASAP7_75t_R   g0614( .A (n1011), .B (n1015), .Y (n1017) );
  INVx1_ASAP7_75t_R      g0615( .A (x57), .Y (n315) );
  XNOR2xp5_ASAP7_75t_R   g0616( .A (n315), .B (x185), .Y (n1022) );
  XNOR2xp5_ASAP7_75t_R   g0617( .A (n1017), .B (n1022), .Y (y57) );
  INVx1_ASAP7_75t_R      g0618( .A (x185), .Y (n443) );
  NOR2xp33_ASAP7_75t_R   g0619( .A (n315), .B (n443), .Y (n1020) );
  NAND2xp33_ASAP7_75t_R  g0620( .A (x56), .B (x184), .Y (n1012) );
  NOR2xp33_ASAP7_75t_R   g0621( .A (x57), .B (x185), .Y (n1018) );
  NAND2xp33_ASAP7_75t_R  g0622( .A (n314), .B (n442), .Y (n1010) );
  OAI21xp33_ASAP7_75t_R  g0623( .A1 (n1002), .A2 (n1006), .B (n1010), .Y (n1016) );
  AOI21xp33_ASAP7_75t_R  g0624( .A1 (n1012), .B (n1018), .A2 (n1016), .Y (n1024) );
  NOR2xp33_ASAP7_75t_R   g0625( .A (n1020), .B (n1024), .Y (n1026) );
  INVx1_ASAP7_75t_R      g0626( .A (x58), .Y (n316) );
  XNOR2xp5_ASAP7_75t_R   g0627( .A (n316), .B (x186), .Y (n1031) );
  XNOR2xp5_ASAP7_75t_R   g0628( .A (n1026), .B (n1031), .Y (y58) );
  INVx1_ASAP7_75t_R      g0629( .A (x186), .Y (n444) );
  NOR2xp33_ASAP7_75t_R   g0630( .A (n316), .B (n444), .Y (n1029) );
  NAND2xp33_ASAP7_75t_R  g0631( .A (x57), .B (x185), .Y (n1021) );
  NOR2xp33_ASAP7_75t_R   g0632( .A (x58), .B (x186), .Y (n1027) );
  NAND2xp33_ASAP7_75t_R  g0633( .A (n315), .B (n443), .Y (n1019) );
  OAI21xp33_ASAP7_75t_R  g0634( .A1 (n1011), .A2 (n1015), .B (n1019), .Y (n1025) );
  AOI21xp33_ASAP7_75t_R  g0635( .A1 (n1021), .B (n1027), .A2 (n1025), .Y (n1033) );
  NOR2xp33_ASAP7_75t_R   g0636( .A (n1029), .B (n1033), .Y (n1035) );
  INVx1_ASAP7_75t_R      g0637( .A (x59), .Y (n317) );
  XNOR2xp5_ASAP7_75t_R   g0638( .A (n317), .B (x187), .Y (n1040) );
  XNOR2xp5_ASAP7_75t_R   g0639( .A (n1035), .B (n1040), .Y (y59) );
  INVx1_ASAP7_75t_R      g0640( .A (x187), .Y (n445) );
  NOR2xp33_ASAP7_75t_R   g0641( .A (n317), .B (n445), .Y (n1038) );
  NAND2xp33_ASAP7_75t_R  g0642( .A (x58), .B (x186), .Y (n1030) );
  NOR2xp33_ASAP7_75t_R   g0643( .A (x59), .B (x187), .Y (n1036) );
  NAND2xp33_ASAP7_75t_R  g0644( .A (n316), .B (n444), .Y (n1028) );
  OAI21xp33_ASAP7_75t_R  g0645( .A1 (n1020), .A2 (n1024), .B (n1028), .Y (n1034) );
  AOI21xp33_ASAP7_75t_R  g0646( .A1 (n1030), .B (n1036), .A2 (n1034), .Y (n1042) );
  NOR2xp33_ASAP7_75t_R   g0647( .A (n1038), .B (n1042), .Y (n1044) );
  INVx1_ASAP7_75t_R      g0648( .A (x60), .Y (n318) );
  XNOR2xp5_ASAP7_75t_R   g0649( .A (n318), .B (x188), .Y (n1049) );
  XNOR2xp5_ASAP7_75t_R   g0650( .A (n1044), .B (n1049), .Y (y60) );
  INVx1_ASAP7_75t_R      g0651( .A (x188), .Y (n446) );
  NOR2xp33_ASAP7_75t_R   g0652( .A (n318), .B (n446), .Y (n1047) );
  NAND2xp33_ASAP7_75t_R  g0653( .A (x59), .B (x187), .Y (n1039) );
  NOR2xp33_ASAP7_75t_R   g0654( .A (x60), .B (x188), .Y (n1045) );
  NAND2xp33_ASAP7_75t_R  g0655( .A (n317), .B (n445), .Y (n1037) );
  OAI21xp33_ASAP7_75t_R  g0656( .A1 (n1029), .A2 (n1033), .B (n1037), .Y (n1043) );
  AOI21xp33_ASAP7_75t_R  g0657( .A1 (n1039), .B (n1045), .A2 (n1043), .Y (n1051) );
  NOR2xp33_ASAP7_75t_R   g0658( .A (n1047), .B (n1051), .Y (n1053) );
  INVx1_ASAP7_75t_R      g0659( .A (x61), .Y (n319) );
  XNOR2xp5_ASAP7_75t_R   g0660( .A (n319), .B (x189), .Y (n1058) );
  XNOR2xp5_ASAP7_75t_R   g0661( .A (n1053), .B (n1058), .Y (y61) );
  INVx1_ASAP7_75t_R      g0662( .A (x189), .Y (n447) );
  NOR2xp33_ASAP7_75t_R   g0663( .A (n319), .B (n447), .Y (n1056) );
  NAND2xp33_ASAP7_75t_R  g0664( .A (x60), .B (x188), .Y (n1048) );
  NOR2xp33_ASAP7_75t_R   g0665( .A (x61), .B (x189), .Y (n1054) );
  NAND2xp33_ASAP7_75t_R  g0666( .A (n318), .B (n446), .Y (n1046) );
  OAI21xp33_ASAP7_75t_R  g0667( .A1 (n1038), .A2 (n1042), .B (n1046), .Y (n1052) );
  AOI21xp33_ASAP7_75t_R  g0668( .A1 (n1048), .B (n1054), .A2 (n1052), .Y (n1060) );
  NOR2xp33_ASAP7_75t_R   g0669( .A (n1056), .B (n1060), .Y (n1062) );
  INVx1_ASAP7_75t_R      g0670( .A (x62), .Y (n320) );
  XNOR2xp5_ASAP7_75t_R   g0671( .A (n320), .B (x190), .Y (n1067) );
  XNOR2xp5_ASAP7_75t_R   g0672( .A (n1062), .B (n1067), .Y (y62) );
  INVx1_ASAP7_75t_R      g0673( .A (x190), .Y (n448) );
  NOR2xp33_ASAP7_75t_R   g0674( .A (n320), .B (n448), .Y (n1065) );
  NAND2xp33_ASAP7_75t_R  g0675( .A (x61), .B (x189), .Y (n1057) );
  NOR2xp33_ASAP7_75t_R   g0676( .A (x62), .B (x190), .Y (n1063) );
  NAND2xp33_ASAP7_75t_R  g0677( .A (n319), .B (n447), .Y (n1055) );
  OAI21xp33_ASAP7_75t_R  g0678( .A1 (n1047), .A2 (n1051), .B (n1055), .Y (n1061) );
  AOI21xp33_ASAP7_75t_R  g0679( .A1 (n1057), .B (n1063), .A2 (n1061), .Y (n1069) );
  NOR2xp33_ASAP7_75t_R   g0680( .A (n1065), .B (n1069), .Y (n1071) );
  INVx1_ASAP7_75t_R      g0681( .A (x63), .Y (n321) );
  XNOR2xp5_ASAP7_75t_R   g0682( .A (n321), .B (x191), .Y (n1076) );
  XNOR2xp5_ASAP7_75t_R   g0683( .A (n1071), .B (n1076), .Y (y63) );
  INVx1_ASAP7_75t_R      g0684( .A (x191), .Y (n449) );
  NOR2xp33_ASAP7_75t_R   g0685( .A (n321), .B (n449), .Y (n1074) );
  NAND2xp33_ASAP7_75t_R  g0686( .A (x62), .B (x190), .Y (n1066) );
  NOR2xp33_ASAP7_75t_R   g0687( .A (x63), .B (x191), .Y (n1072) );
  NAND2xp33_ASAP7_75t_R  g0688( .A (n320), .B (n448), .Y (n1064) );
  OAI21xp33_ASAP7_75t_R  g0689( .A1 (n1056), .A2 (n1060), .B (n1064), .Y (n1070) );
  AOI21xp33_ASAP7_75t_R  g0690( .A1 (n1066), .B (n1072), .A2 (n1070), .Y (n1078) );
  NOR2xp33_ASAP7_75t_R   g0691( .A (n1074), .B (n1078), .Y (n1080) );
  INVx1_ASAP7_75t_R      g0692( .A (x64), .Y (n322) );
  XNOR2xp5_ASAP7_75t_R   g0693( .A (n322), .B (x192), .Y (n1085) );
  XNOR2xp5_ASAP7_75t_R   g0694( .A (n1080), .B (n1085), .Y (y64) );
  INVx1_ASAP7_75t_R      g0695( .A (x192), .Y (n450) );
  NOR2xp33_ASAP7_75t_R   g0696( .A (n322), .B (n450), .Y (n1083) );
  NAND2xp33_ASAP7_75t_R  g0697( .A (x63), .B (x191), .Y (n1075) );
  NOR2xp33_ASAP7_75t_R   g0698( .A (x64), .B (x192), .Y (n1081) );
  NAND2xp33_ASAP7_75t_R  g0699( .A (n321), .B (n449), .Y (n1073) );
  OAI21xp33_ASAP7_75t_R  g0700( .A1 (n1065), .A2 (n1069), .B (n1073), .Y (n1079) );
  AOI21xp33_ASAP7_75t_R  g0701( .A1 (n1075), .B (n1081), .A2 (n1079), .Y (n1087) );
  NOR2xp33_ASAP7_75t_R   g0702( .A (n1083), .B (n1087), .Y (n1089) );
  INVx1_ASAP7_75t_R      g0703( .A (x65), .Y (n323) );
  XNOR2xp5_ASAP7_75t_R   g0704( .A (n323), .B (x193), .Y (n1094) );
  XNOR2xp5_ASAP7_75t_R   g0705( .A (n1089), .B (n1094), .Y (y65) );
  INVx1_ASAP7_75t_R      g0706( .A (x193), .Y (n451) );
  NOR2xp33_ASAP7_75t_R   g0707( .A (n323), .B (n451), .Y (n1092) );
  NAND2xp33_ASAP7_75t_R  g0708( .A (x64), .B (x192), .Y (n1084) );
  NOR2xp33_ASAP7_75t_R   g0709( .A (x65), .B (x193), .Y (n1090) );
  NAND2xp33_ASAP7_75t_R  g0710( .A (n322), .B (n450), .Y (n1082) );
  OAI21xp33_ASAP7_75t_R  g0711( .A1 (n1074), .A2 (n1078), .B (n1082), .Y (n1088) );
  AOI21xp33_ASAP7_75t_R  g0712( .A1 (n1084), .B (n1090), .A2 (n1088), .Y (n1096) );
  NOR2xp33_ASAP7_75t_R   g0713( .A (n1092), .B (n1096), .Y (n1098) );
  INVx1_ASAP7_75t_R      g0714( .A (x66), .Y (n324) );
  XNOR2xp5_ASAP7_75t_R   g0715( .A (n324), .B (x194), .Y (n1103) );
  XNOR2xp5_ASAP7_75t_R   g0716( .A (n1098), .B (n1103), .Y (y66) );
  INVx1_ASAP7_75t_R      g0717( .A (x194), .Y (n452) );
  NOR2xp33_ASAP7_75t_R   g0718( .A (n324), .B (n452), .Y (n1101) );
  NAND2xp33_ASAP7_75t_R  g0719( .A (x65), .B (x193), .Y (n1093) );
  NOR2xp33_ASAP7_75t_R   g0720( .A (x66), .B (x194), .Y (n1099) );
  NAND2xp33_ASAP7_75t_R  g0721( .A (n323), .B (n451), .Y (n1091) );
  OAI21xp33_ASAP7_75t_R  g0722( .A1 (n1083), .A2 (n1087), .B (n1091), .Y (n1097) );
  AOI21xp33_ASAP7_75t_R  g0723( .A1 (n1093), .B (n1099), .A2 (n1097), .Y (n1105) );
  NOR2xp33_ASAP7_75t_R   g0724( .A (n1101), .B (n1105), .Y (n1107) );
  INVx1_ASAP7_75t_R      g0725( .A (x67), .Y (n325) );
  XNOR2xp5_ASAP7_75t_R   g0726( .A (n325), .B (x195), .Y (n1112) );
  XNOR2xp5_ASAP7_75t_R   g0727( .A (n1107), .B (n1112), .Y (y67) );
  INVx1_ASAP7_75t_R      g0728( .A (x195), .Y (n453) );
  NOR2xp33_ASAP7_75t_R   g0729( .A (n325), .B (n453), .Y (n1110) );
  NAND2xp33_ASAP7_75t_R  g0730( .A (x66), .B (x194), .Y (n1102) );
  NOR2xp33_ASAP7_75t_R   g0731( .A (x67), .B (x195), .Y (n1108) );
  NAND2xp33_ASAP7_75t_R  g0732( .A (n324), .B (n452), .Y (n1100) );
  OAI21xp33_ASAP7_75t_R  g0733( .A1 (n1092), .A2 (n1096), .B (n1100), .Y (n1106) );
  AOI21xp33_ASAP7_75t_R  g0734( .A1 (n1102), .B (n1108), .A2 (n1106), .Y (n1114) );
  NOR2xp33_ASAP7_75t_R   g0735( .A (n1110), .B (n1114), .Y (n1116) );
  INVx1_ASAP7_75t_R      g0736( .A (x68), .Y (n326) );
  XNOR2xp5_ASAP7_75t_R   g0737( .A (n326), .B (x196), .Y (n1121) );
  XNOR2xp5_ASAP7_75t_R   g0738( .A (n1116), .B (n1121), .Y (y68) );
  INVx1_ASAP7_75t_R      g0739( .A (x196), .Y (n454) );
  NOR2xp33_ASAP7_75t_R   g0740( .A (n326), .B (n454), .Y (n1119) );
  NAND2xp33_ASAP7_75t_R  g0741( .A (x67), .B (x195), .Y (n1111) );
  NOR2xp33_ASAP7_75t_R   g0742( .A (x68), .B (x196), .Y (n1117) );
  NAND2xp33_ASAP7_75t_R  g0743( .A (n325), .B (n453), .Y (n1109) );
  OAI21xp33_ASAP7_75t_R  g0744( .A1 (n1101), .A2 (n1105), .B (n1109), .Y (n1115) );
  AOI21xp33_ASAP7_75t_R  g0745( .A1 (n1111), .B (n1117), .A2 (n1115), .Y (n1123) );
  NOR2xp33_ASAP7_75t_R   g0746( .A (n1119), .B (n1123), .Y (n1125) );
  INVx1_ASAP7_75t_R      g0747( .A (x69), .Y (n327) );
  XNOR2xp5_ASAP7_75t_R   g0748( .A (n327), .B (x197), .Y (n1130) );
  XNOR2xp5_ASAP7_75t_R   g0749( .A (n1125), .B (n1130), .Y (y69) );
  INVx1_ASAP7_75t_R      g0750( .A (x197), .Y (n455) );
  NOR2xp33_ASAP7_75t_R   g0751( .A (n327), .B (n455), .Y (n1128) );
  NAND2xp33_ASAP7_75t_R  g0752( .A (x68), .B (x196), .Y (n1120) );
  NOR2xp33_ASAP7_75t_R   g0753( .A (x69), .B (x197), .Y (n1126) );
  NAND2xp33_ASAP7_75t_R  g0754( .A (n326), .B (n454), .Y (n1118) );
  OAI21xp33_ASAP7_75t_R  g0755( .A1 (n1110), .A2 (n1114), .B (n1118), .Y (n1124) );
  AOI21xp33_ASAP7_75t_R  g0756( .A1 (n1120), .B (n1126), .A2 (n1124), .Y (n1132) );
  NOR2xp33_ASAP7_75t_R   g0757( .A (n1128), .B (n1132), .Y (n1134) );
  INVx1_ASAP7_75t_R      g0758( .A (x70), .Y (n328) );
  XNOR2xp5_ASAP7_75t_R   g0759( .A (n328), .B (x198), .Y (n1139) );
  XNOR2xp5_ASAP7_75t_R   g0760( .A (n1134), .B (n1139), .Y (y70) );
  INVx1_ASAP7_75t_R      g0761( .A (x198), .Y (n456) );
  NOR2xp33_ASAP7_75t_R   g0762( .A (n328), .B (n456), .Y (n1137) );
  NAND2xp33_ASAP7_75t_R  g0763( .A (x69), .B (x197), .Y (n1129) );
  NOR2xp33_ASAP7_75t_R   g0764( .A (x70), .B (x198), .Y (n1135) );
  NAND2xp33_ASAP7_75t_R  g0765( .A (n327), .B (n455), .Y (n1127) );
  OAI21xp33_ASAP7_75t_R  g0766( .A1 (n1119), .A2 (n1123), .B (n1127), .Y (n1133) );
  AOI21xp33_ASAP7_75t_R  g0767( .A1 (n1129), .B (n1135), .A2 (n1133), .Y (n1141) );
  NOR2xp33_ASAP7_75t_R   g0768( .A (n1137), .B (n1141), .Y (n1143) );
  INVx1_ASAP7_75t_R      g0769( .A (x71), .Y (n329) );
  XNOR2xp5_ASAP7_75t_R   g0770( .A (n329), .B (x199), .Y (n1148) );
  XNOR2xp5_ASAP7_75t_R   g0771( .A (n1143), .B (n1148), .Y (y71) );
  INVx1_ASAP7_75t_R      g0772( .A (x199), .Y (n457) );
  NOR2xp33_ASAP7_75t_R   g0773( .A (n329), .B (n457), .Y (n1146) );
  NAND2xp33_ASAP7_75t_R  g0774( .A (x70), .B (x198), .Y (n1138) );
  NOR2xp33_ASAP7_75t_R   g0775( .A (x71), .B (x199), .Y (n1144) );
  NAND2xp33_ASAP7_75t_R  g0776( .A (n328), .B (n456), .Y (n1136) );
  OAI21xp33_ASAP7_75t_R  g0777( .A1 (n1128), .A2 (n1132), .B (n1136), .Y (n1142) );
  AOI21xp33_ASAP7_75t_R  g0778( .A1 (n1138), .B (n1144), .A2 (n1142), .Y (n1150) );
  NOR2xp33_ASAP7_75t_R   g0779( .A (n1146), .B (n1150), .Y (n1152) );
  INVx1_ASAP7_75t_R      g0780( .A (x72), .Y (n330) );
  XNOR2xp5_ASAP7_75t_R   g0781( .A (n330), .B (x200), .Y (n1157) );
  XNOR2xp5_ASAP7_75t_R   g0782( .A (n1152), .B (n1157), .Y (y72) );
  INVx1_ASAP7_75t_R      g0783( .A (x200), .Y (n458) );
  NOR2xp33_ASAP7_75t_R   g0784( .A (n330), .B (n458), .Y (n1155) );
  NAND2xp33_ASAP7_75t_R  g0785( .A (x71), .B (x199), .Y (n1147) );
  NOR2xp33_ASAP7_75t_R   g0786( .A (x72), .B (x200), .Y (n1153) );
  NAND2xp33_ASAP7_75t_R  g0787( .A (n329), .B (n457), .Y (n1145) );
  OAI21xp33_ASAP7_75t_R  g0788( .A1 (n1137), .A2 (n1141), .B (n1145), .Y (n1151) );
  AOI21xp33_ASAP7_75t_R  g0789( .A1 (n1147), .B (n1153), .A2 (n1151), .Y (n1159) );
  NOR2xp33_ASAP7_75t_R   g0790( .A (n1155), .B (n1159), .Y (n1161) );
  INVx1_ASAP7_75t_R      g0791( .A (x73), .Y (n331) );
  XNOR2xp5_ASAP7_75t_R   g0792( .A (n331), .B (x201), .Y (n1166) );
  XNOR2xp5_ASAP7_75t_R   g0793( .A (n1161), .B (n1166), .Y (y73) );
  INVx1_ASAP7_75t_R      g0794( .A (x201), .Y (n459) );
  NOR2xp33_ASAP7_75t_R   g0795( .A (n331), .B (n459), .Y (n1164) );
  NAND2xp33_ASAP7_75t_R  g0796( .A (x72), .B (x200), .Y (n1156) );
  NOR2xp33_ASAP7_75t_R   g0797( .A (x73), .B (x201), .Y (n1162) );
  NAND2xp33_ASAP7_75t_R  g0798( .A (n330), .B (n458), .Y (n1154) );
  OAI21xp33_ASAP7_75t_R  g0799( .A1 (n1146), .A2 (n1150), .B (n1154), .Y (n1160) );
  AOI21xp33_ASAP7_75t_R  g0800( .A1 (n1156), .B (n1162), .A2 (n1160), .Y (n1168) );
  NOR2xp33_ASAP7_75t_R   g0801( .A (n1164), .B (n1168), .Y (n1170) );
  INVx1_ASAP7_75t_R      g0802( .A (x74), .Y (n332) );
  XNOR2xp5_ASAP7_75t_R   g0803( .A (n332), .B (x202), .Y (n1175) );
  XNOR2xp5_ASAP7_75t_R   g0804( .A (n1170), .B (n1175), .Y (y74) );
  INVx1_ASAP7_75t_R      g0805( .A (x202), .Y (n460) );
  NOR2xp33_ASAP7_75t_R   g0806( .A (n332), .B (n460), .Y (n1173) );
  NAND2xp33_ASAP7_75t_R  g0807( .A (x73), .B (x201), .Y (n1165) );
  NOR2xp33_ASAP7_75t_R   g0808( .A (x74), .B (x202), .Y (n1171) );
  NAND2xp33_ASAP7_75t_R  g0809( .A (n331), .B (n459), .Y (n1163) );
  OAI21xp33_ASAP7_75t_R  g0810( .A1 (n1155), .A2 (n1159), .B (n1163), .Y (n1169) );
  AOI21xp33_ASAP7_75t_R  g0811( .A1 (n1165), .B (n1171), .A2 (n1169), .Y (n1177) );
  NOR2xp33_ASAP7_75t_R   g0812( .A (n1173), .B (n1177), .Y (n1179) );
  INVx1_ASAP7_75t_R      g0813( .A (x75), .Y (n333) );
  XNOR2xp5_ASAP7_75t_R   g0814( .A (n333), .B (x203), .Y (n1184) );
  XNOR2xp5_ASAP7_75t_R   g0815( .A (n1179), .B (n1184), .Y (y75) );
  INVx1_ASAP7_75t_R      g0816( .A (x203), .Y (n461) );
  NOR2xp33_ASAP7_75t_R   g0817( .A (n333), .B (n461), .Y (n1182) );
  NAND2xp33_ASAP7_75t_R  g0818( .A (x74), .B (x202), .Y (n1174) );
  NOR2xp33_ASAP7_75t_R   g0819( .A (x75), .B (x203), .Y (n1180) );
  NAND2xp33_ASAP7_75t_R  g0820( .A (n332), .B (n460), .Y (n1172) );
  OAI21xp33_ASAP7_75t_R  g0821( .A1 (n1164), .A2 (n1168), .B (n1172), .Y (n1178) );
  AOI21xp33_ASAP7_75t_R  g0822( .A1 (n1174), .B (n1180), .A2 (n1178), .Y (n1186) );
  NOR2xp33_ASAP7_75t_R   g0823( .A (n1182), .B (n1186), .Y (n1188) );
  INVx1_ASAP7_75t_R      g0824( .A (x76), .Y (n334) );
  XNOR2xp5_ASAP7_75t_R   g0825( .A (n334), .B (x204), .Y (n1193) );
  XNOR2xp5_ASAP7_75t_R   g0826( .A (n1188), .B (n1193), .Y (y76) );
  INVx1_ASAP7_75t_R      g0827( .A (x204), .Y (n462) );
  NOR2xp33_ASAP7_75t_R   g0828( .A (n334), .B (n462), .Y (n1191) );
  NAND2xp33_ASAP7_75t_R  g0829( .A (x75), .B (x203), .Y (n1183) );
  NOR2xp33_ASAP7_75t_R   g0830( .A (x76), .B (x204), .Y (n1189) );
  NAND2xp33_ASAP7_75t_R  g0831( .A (n333), .B (n461), .Y (n1181) );
  OAI21xp33_ASAP7_75t_R  g0832( .A1 (n1173), .A2 (n1177), .B (n1181), .Y (n1187) );
  AOI21xp33_ASAP7_75t_R  g0833( .A1 (n1183), .B (n1189), .A2 (n1187), .Y (n1195) );
  NOR2xp33_ASAP7_75t_R   g0834( .A (n1191), .B (n1195), .Y (n1197) );
  INVx1_ASAP7_75t_R      g0835( .A (x77), .Y (n335) );
  XNOR2xp5_ASAP7_75t_R   g0836( .A (n335), .B (x205), .Y (n1202) );
  XNOR2xp5_ASAP7_75t_R   g0837( .A (n1197), .B (n1202), .Y (y77) );
  INVx1_ASAP7_75t_R      g0838( .A (x205), .Y (n463) );
  NOR2xp33_ASAP7_75t_R   g0839( .A (n335), .B (n463), .Y (n1200) );
  NAND2xp33_ASAP7_75t_R  g0840( .A (x76), .B (x204), .Y (n1192) );
  NOR2xp33_ASAP7_75t_R   g0841( .A (x77), .B (x205), .Y (n1198) );
  NAND2xp33_ASAP7_75t_R  g0842( .A (n334), .B (n462), .Y (n1190) );
  OAI21xp33_ASAP7_75t_R  g0843( .A1 (n1182), .A2 (n1186), .B (n1190), .Y (n1196) );
  AOI21xp33_ASAP7_75t_R  g0844( .A1 (n1192), .B (n1198), .A2 (n1196), .Y (n1204) );
  NOR2xp33_ASAP7_75t_R   g0845( .A (n1200), .B (n1204), .Y (n1206) );
  INVx1_ASAP7_75t_R      g0846( .A (x78), .Y (n336) );
  XNOR2xp5_ASAP7_75t_R   g0847( .A (n336), .B (x206), .Y (n1211) );
  XNOR2xp5_ASAP7_75t_R   g0848( .A (n1206), .B (n1211), .Y (y78) );
  INVx1_ASAP7_75t_R      g0849( .A (x206), .Y (n464) );
  NOR2xp33_ASAP7_75t_R   g0850( .A (n336), .B (n464), .Y (n1209) );
  NAND2xp33_ASAP7_75t_R  g0851( .A (x77), .B (x205), .Y (n1201) );
  NOR2xp33_ASAP7_75t_R   g0852( .A (x78), .B (x206), .Y (n1207) );
  NAND2xp33_ASAP7_75t_R  g0853( .A (n335), .B (n463), .Y (n1199) );
  OAI21xp33_ASAP7_75t_R  g0854( .A1 (n1191), .A2 (n1195), .B (n1199), .Y (n1205) );
  AOI21xp33_ASAP7_75t_R  g0855( .A1 (n1201), .B (n1207), .A2 (n1205), .Y (n1213) );
  NOR2xp33_ASAP7_75t_R   g0856( .A (n1209), .B (n1213), .Y (n1215) );
  INVx1_ASAP7_75t_R      g0857( .A (x79), .Y (n337) );
  XNOR2xp5_ASAP7_75t_R   g0858( .A (n337), .B (x207), .Y (n1220) );
  XNOR2xp5_ASAP7_75t_R   g0859( .A (n1215), .B (n1220), .Y (y79) );
  INVx1_ASAP7_75t_R      g0860( .A (x207), .Y (n465) );
  NOR2xp33_ASAP7_75t_R   g0861( .A (n337), .B (n465), .Y (n1218) );
  NAND2xp33_ASAP7_75t_R  g0862( .A (x78), .B (x206), .Y (n1210) );
  NOR2xp33_ASAP7_75t_R   g0863( .A (x79), .B (x207), .Y (n1216) );
  NAND2xp33_ASAP7_75t_R  g0864( .A (n336), .B (n464), .Y (n1208) );
  OAI21xp33_ASAP7_75t_R  g0865( .A1 (n1200), .A2 (n1204), .B (n1208), .Y (n1214) );
  AOI21xp33_ASAP7_75t_R  g0866( .A1 (n1210), .B (n1216), .A2 (n1214), .Y (n1222) );
  NOR2xp33_ASAP7_75t_R   g0867( .A (n1218), .B (n1222), .Y (n1224) );
  INVx1_ASAP7_75t_R      g0868( .A (x80), .Y (n338) );
  XNOR2xp5_ASAP7_75t_R   g0869( .A (n338), .B (x208), .Y (n1229) );
  XNOR2xp5_ASAP7_75t_R   g0870( .A (n1224), .B (n1229), .Y (y80) );
  INVx1_ASAP7_75t_R      g0871( .A (x208), .Y (n466) );
  NOR2xp33_ASAP7_75t_R   g0872( .A (n338), .B (n466), .Y (n1227) );
  NAND2xp33_ASAP7_75t_R  g0873( .A (x79), .B (x207), .Y (n1219) );
  NOR2xp33_ASAP7_75t_R   g0874( .A (x80), .B (x208), .Y (n1225) );
  NAND2xp33_ASAP7_75t_R  g0875( .A (n337), .B (n465), .Y (n1217) );
  OAI21xp33_ASAP7_75t_R  g0876( .A1 (n1209), .A2 (n1213), .B (n1217), .Y (n1223) );
  AOI21xp33_ASAP7_75t_R  g0877( .A1 (n1219), .B (n1225), .A2 (n1223), .Y (n1231) );
  NOR2xp33_ASAP7_75t_R   g0878( .A (n1227), .B (n1231), .Y (n1233) );
  INVx1_ASAP7_75t_R      g0879( .A (x81), .Y (n339) );
  XNOR2xp5_ASAP7_75t_R   g0880( .A (n339), .B (x209), .Y (n1238) );
  XNOR2xp5_ASAP7_75t_R   g0881( .A (n1233), .B (n1238), .Y (y81) );
  INVx1_ASAP7_75t_R      g0882( .A (x209), .Y (n467) );
  NOR2xp33_ASAP7_75t_R   g0883( .A (n339), .B (n467), .Y (n1236) );
  NAND2xp33_ASAP7_75t_R  g0884( .A (x80), .B (x208), .Y (n1228) );
  NOR2xp33_ASAP7_75t_R   g0885( .A (x81), .B (x209), .Y (n1234) );
  NAND2xp33_ASAP7_75t_R  g0886( .A (n338), .B (n466), .Y (n1226) );
  OAI21xp33_ASAP7_75t_R  g0887( .A1 (n1218), .A2 (n1222), .B (n1226), .Y (n1232) );
  AOI21xp33_ASAP7_75t_R  g0888( .A1 (n1228), .B (n1234), .A2 (n1232), .Y (n1240) );
  NOR2xp33_ASAP7_75t_R   g0889( .A (n1236), .B (n1240), .Y (n1242) );
  INVx1_ASAP7_75t_R      g0890( .A (x82), .Y (n340) );
  XNOR2xp5_ASAP7_75t_R   g0891( .A (n340), .B (x210), .Y (n1247) );
  XNOR2xp5_ASAP7_75t_R   g0892( .A (n1242), .B (n1247), .Y (y82) );
  INVx1_ASAP7_75t_R      g0893( .A (x210), .Y (n468) );
  NOR2xp33_ASAP7_75t_R   g0894( .A (n340), .B (n468), .Y (n1245) );
  NAND2xp33_ASAP7_75t_R  g0895( .A (x81), .B (x209), .Y (n1237) );
  NOR2xp33_ASAP7_75t_R   g0896( .A (x82), .B (x210), .Y (n1243) );
  NAND2xp33_ASAP7_75t_R  g0897( .A (n339), .B (n467), .Y (n1235) );
  OAI21xp33_ASAP7_75t_R  g0898( .A1 (n1227), .A2 (n1231), .B (n1235), .Y (n1241) );
  AOI21xp33_ASAP7_75t_R  g0899( .A1 (n1237), .B (n1243), .A2 (n1241), .Y (n1249) );
  NOR2xp33_ASAP7_75t_R   g0900( .A (n1245), .B (n1249), .Y (n1251) );
  INVx1_ASAP7_75t_R      g0901( .A (x83), .Y (n341) );
  XNOR2xp5_ASAP7_75t_R   g0902( .A (n341), .B (x211), .Y (n1256) );
  XNOR2xp5_ASAP7_75t_R   g0903( .A (n1251), .B (n1256), .Y (y83) );
  INVx1_ASAP7_75t_R      g0904( .A (x211), .Y (n469) );
  NOR2xp33_ASAP7_75t_R   g0905( .A (n341), .B (n469), .Y (n1254) );
  NAND2xp33_ASAP7_75t_R  g0906( .A (x82), .B (x210), .Y (n1246) );
  NOR2xp33_ASAP7_75t_R   g0907( .A (x83), .B (x211), .Y (n1252) );
  NAND2xp33_ASAP7_75t_R  g0908( .A (n340), .B (n468), .Y (n1244) );
  OAI21xp33_ASAP7_75t_R  g0909( .A1 (n1236), .A2 (n1240), .B (n1244), .Y (n1250) );
  AOI21xp33_ASAP7_75t_R  g0910( .A1 (n1246), .B (n1252), .A2 (n1250), .Y (n1258) );
  NOR2xp33_ASAP7_75t_R   g0911( .A (n1254), .B (n1258), .Y (n1260) );
  INVx1_ASAP7_75t_R      g0912( .A (x84), .Y (n342) );
  XNOR2xp5_ASAP7_75t_R   g0913( .A (n342), .B (x212), .Y (n1265) );
  XNOR2xp5_ASAP7_75t_R   g0914( .A (n1260), .B (n1265), .Y (y84) );
  INVx1_ASAP7_75t_R      g0915( .A (x212), .Y (n470) );
  NOR2xp33_ASAP7_75t_R   g0916( .A (n342), .B (n470), .Y (n1263) );
  NAND2xp33_ASAP7_75t_R  g0917( .A (x83), .B (x211), .Y (n1255) );
  NOR2xp33_ASAP7_75t_R   g0918( .A (x84), .B (x212), .Y (n1261) );
  NAND2xp33_ASAP7_75t_R  g0919( .A (n341), .B (n469), .Y (n1253) );
  OAI21xp33_ASAP7_75t_R  g0920( .A1 (n1245), .A2 (n1249), .B (n1253), .Y (n1259) );
  AOI21xp33_ASAP7_75t_R  g0921( .A1 (n1255), .B (n1261), .A2 (n1259), .Y (n1267) );
  NOR2xp33_ASAP7_75t_R   g0922( .A (n1263), .B (n1267), .Y (n1269) );
  INVx1_ASAP7_75t_R      g0923( .A (x85), .Y (n343) );
  XNOR2xp5_ASAP7_75t_R   g0924( .A (n343), .B (x213), .Y (n1274) );
  XNOR2xp5_ASAP7_75t_R   g0925( .A (n1269), .B (n1274), .Y (y85) );
  INVx1_ASAP7_75t_R      g0926( .A (x213), .Y (n471) );
  NOR2xp33_ASAP7_75t_R   g0927( .A (n343), .B (n471), .Y (n1272) );
  NAND2xp33_ASAP7_75t_R  g0928( .A (x84), .B (x212), .Y (n1264) );
  NOR2xp33_ASAP7_75t_R   g0929( .A (x85), .B (x213), .Y (n1270) );
  NAND2xp33_ASAP7_75t_R  g0930( .A (n342), .B (n470), .Y (n1262) );
  OAI21xp33_ASAP7_75t_R  g0931( .A1 (n1254), .A2 (n1258), .B (n1262), .Y (n1268) );
  AOI21xp33_ASAP7_75t_R  g0932( .A1 (n1264), .B (n1270), .A2 (n1268), .Y (n1276) );
  NOR2xp33_ASAP7_75t_R   g0933( .A (n1272), .B (n1276), .Y (n1278) );
  INVx1_ASAP7_75t_R      g0934( .A (x86), .Y (n344) );
  XNOR2xp5_ASAP7_75t_R   g0935( .A (n344), .B (x214), .Y (n1283) );
  XNOR2xp5_ASAP7_75t_R   g0936( .A (n1278), .B (n1283), .Y (y86) );
  INVx1_ASAP7_75t_R      g0937( .A (x214), .Y (n472) );
  NOR2xp33_ASAP7_75t_R   g0938( .A (n344), .B (n472), .Y (n1281) );
  NAND2xp33_ASAP7_75t_R  g0939( .A (x85), .B (x213), .Y (n1273) );
  NOR2xp33_ASAP7_75t_R   g0940( .A (x86), .B (x214), .Y (n1279) );
  NAND2xp33_ASAP7_75t_R  g0941( .A (n343), .B (n471), .Y (n1271) );
  OAI21xp33_ASAP7_75t_R  g0942( .A1 (n1263), .A2 (n1267), .B (n1271), .Y (n1277) );
  AOI21xp33_ASAP7_75t_R  g0943( .A1 (n1273), .B (n1279), .A2 (n1277), .Y (n1285) );
  NOR2xp33_ASAP7_75t_R   g0944( .A (n1281), .B (n1285), .Y (n1287) );
  INVx1_ASAP7_75t_R      g0945( .A (x87), .Y (n345) );
  XNOR2xp5_ASAP7_75t_R   g0946( .A (n345), .B (x215), .Y (n1292) );
  XNOR2xp5_ASAP7_75t_R   g0947( .A (n1287), .B (n1292), .Y (y87) );
  INVx1_ASAP7_75t_R      g0948( .A (x215), .Y (n473) );
  NOR2xp33_ASAP7_75t_R   g0949( .A (n345), .B (n473), .Y (n1290) );
  NAND2xp33_ASAP7_75t_R  g0950( .A (x86), .B (x214), .Y (n1282) );
  NOR2xp33_ASAP7_75t_R   g0951( .A (x87), .B (x215), .Y (n1288) );
  NAND2xp33_ASAP7_75t_R  g0952( .A (n344), .B (n472), .Y (n1280) );
  OAI21xp33_ASAP7_75t_R  g0953( .A1 (n1272), .A2 (n1276), .B (n1280), .Y (n1286) );
  AOI21xp33_ASAP7_75t_R  g0954( .A1 (n1282), .B (n1288), .A2 (n1286), .Y (n1294) );
  NOR2xp33_ASAP7_75t_R   g0955( .A (n1290), .B (n1294), .Y (n1296) );
  INVx1_ASAP7_75t_R      g0956( .A (x88), .Y (n346) );
  XNOR2xp5_ASAP7_75t_R   g0957( .A (n346), .B (x216), .Y (n1301) );
  XNOR2xp5_ASAP7_75t_R   g0958( .A (n1296), .B (n1301), .Y (y88) );
  INVx1_ASAP7_75t_R      g0959( .A (x216), .Y (n474) );
  NOR2xp33_ASAP7_75t_R   g0960( .A (n346), .B (n474), .Y (n1299) );
  NAND2xp33_ASAP7_75t_R  g0961( .A (x87), .B (x215), .Y (n1291) );
  NOR2xp33_ASAP7_75t_R   g0962( .A (x88), .B (x216), .Y (n1297) );
  NAND2xp33_ASAP7_75t_R  g0963( .A (n345), .B (n473), .Y (n1289) );
  OAI21xp33_ASAP7_75t_R  g0964( .A1 (n1281), .A2 (n1285), .B (n1289), .Y (n1295) );
  AOI21xp33_ASAP7_75t_R  g0965( .A1 (n1291), .B (n1297), .A2 (n1295), .Y (n1303) );
  NOR2xp33_ASAP7_75t_R   g0966( .A (n1299), .B (n1303), .Y (n1305) );
  INVx1_ASAP7_75t_R      g0967( .A (x89), .Y (n347) );
  XNOR2xp5_ASAP7_75t_R   g0968( .A (n347), .B (x217), .Y (n1310) );
  XNOR2xp5_ASAP7_75t_R   g0969( .A (n1305), .B (n1310), .Y (y89) );
  INVx1_ASAP7_75t_R      g0970( .A (x217), .Y (n475) );
  NOR2xp33_ASAP7_75t_R   g0971( .A (n347), .B (n475), .Y (n1308) );
  NAND2xp33_ASAP7_75t_R  g0972( .A (x88), .B (x216), .Y (n1300) );
  NOR2xp33_ASAP7_75t_R   g0973( .A (x89), .B (x217), .Y (n1306) );
  NAND2xp33_ASAP7_75t_R  g0974( .A (n346), .B (n474), .Y (n1298) );
  OAI21xp33_ASAP7_75t_R  g0975( .A1 (n1290), .A2 (n1294), .B (n1298), .Y (n1304) );
  AOI21xp33_ASAP7_75t_R  g0976( .A1 (n1300), .B (n1306), .A2 (n1304), .Y (n1312) );
  NOR2xp33_ASAP7_75t_R   g0977( .A (n1308), .B (n1312), .Y (n1314) );
  INVx1_ASAP7_75t_R      g0978( .A (x90), .Y (n348) );
  XNOR2xp5_ASAP7_75t_R   g0979( .A (n348), .B (x218), .Y (n1319) );
  XNOR2xp5_ASAP7_75t_R   g0980( .A (n1314), .B (n1319), .Y (y90) );
  INVx1_ASAP7_75t_R      g0981( .A (x218), .Y (n476) );
  NOR2xp33_ASAP7_75t_R   g0982( .A (n348), .B (n476), .Y (n1317) );
  NAND2xp33_ASAP7_75t_R  g0983( .A (x89), .B (x217), .Y (n1309) );
  NOR2xp33_ASAP7_75t_R   g0984( .A (x90), .B (x218), .Y (n1315) );
  NAND2xp33_ASAP7_75t_R  g0985( .A (n347), .B (n475), .Y (n1307) );
  OAI21xp33_ASAP7_75t_R  g0986( .A1 (n1299), .A2 (n1303), .B (n1307), .Y (n1313) );
  AOI21xp33_ASAP7_75t_R  g0987( .A1 (n1309), .B (n1315), .A2 (n1313), .Y (n1321) );
  NOR2xp33_ASAP7_75t_R   g0988( .A (n1317), .B (n1321), .Y (n1323) );
  INVx1_ASAP7_75t_R      g0989( .A (x91), .Y (n349) );
  XNOR2xp5_ASAP7_75t_R   g0990( .A (n349), .B (x219), .Y (n1328) );
  XNOR2xp5_ASAP7_75t_R   g0991( .A (n1323), .B (n1328), .Y (y91) );
  INVx1_ASAP7_75t_R      g0992( .A (x219), .Y (n477) );
  NOR2xp33_ASAP7_75t_R   g0993( .A (n349), .B (n477), .Y (n1326) );
  NAND2xp33_ASAP7_75t_R  g0994( .A (x90), .B (x218), .Y (n1318) );
  NOR2xp33_ASAP7_75t_R   g0995( .A (x91), .B (x219), .Y (n1324) );
  NAND2xp33_ASAP7_75t_R  g0996( .A (n348), .B (n476), .Y (n1316) );
  OAI21xp33_ASAP7_75t_R  g0997( .A1 (n1308), .A2 (n1312), .B (n1316), .Y (n1322) );
  AOI21xp33_ASAP7_75t_R  g0998( .A1 (n1318), .B (n1324), .A2 (n1322), .Y (n1330) );
  NOR2xp33_ASAP7_75t_R   g0999( .A (n1326), .B (n1330), .Y (n1332) );
  INVx1_ASAP7_75t_R      g1000( .A (x92), .Y (n350) );
  XNOR2xp5_ASAP7_75t_R   g1001( .A (n350), .B (x220), .Y (n1337) );
  XNOR2xp5_ASAP7_75t_R   g1002( .A (n1332), .B (n1337), .Y (y92) );
  INVx1_ASAP7_75t_R      g1003( .A (x220), .Y (n478) );
  NOR2xp33_ASAP7_75t_R   g1004( .A (n350), .B (n478), .Y (n1335) );
  NAND2xp33_ASAP7_75t_R  g1005( .A (x91), .B (x219), .Y (n1327) );
  NOR2xp33_ASAP7_75t_R   g1006( .A (x92), .B (x220), .Y (n1333) );
  NAND2xp33_ASAP7_75t_R  g1007( .A (n349), .B (n477), .Y (n1325) );
  OAI21xp33_ASAP7_75t_R  g1008( .A1 (n1317), .A2 (n1321), .B (n1325), .Y (n1331) );
  AOI21xp33_ASAP7_75t_R  g1009( .A1 (n1327), .B (n1333), .A2 (n1331), .Y (n1339) );
  NOR2xp33_ASAP7_75t_R   g1010( .A (n1335), .B (n1339), .Y (n1341) );
  INVx1_ASAP7_75t_R      g1011( .A (x93), .Y (n351) );
  XNOR2xp5_ASAP7_75t_R   g1012( .A (n351), .B (x221), .Y (n1346) );
  XNOR2xp5_ASAP7_75t_R   g1013( .A (n1341), .B (n1346), .Y (y93) );
  INVx1_ASAP7_75t_R      g1014( .A (x221), .Y (n479) );
  NOR2xp33_ASAP7_75t_R   g1015( .A (n351), .B (n479), .Y (n1344) );
  NAND2xp33_ASAP7_75t_R  g1016( .A (x92), .B (x220), .Y (n1336) );
  NOR2xp33_ASAP7_75t_R   g1017( .A (x93), .B (x221), .Y (n1342) );
  NAND2xp33_ASAP7_75t_R  g1018( .A (n350), .B (n478), .Y (n1334) );
  OAI21xp33_ASAP7_75t_R  g1019( .A1 (n1326), .A2 (n1330), .B (n1334), .Y (n1340) );
  AOI21xp33_ASAP7_75t_R  g1020( .A1 (n1336), .B (n1342), .A2 (n1340), .Y (n1348) );
  NOR2xp33_ASAP7_75t_R   g1021( .A (n1344), .B (n1348), .Y (n1350) );
  INVx1_ASAP7_75t_R      g1022( .A (x94), .Y (n352) );
  XNOR2xp5_ASAP7_75t_R   g1023( .A (n352), .B (x222), .Y (n1355) );
  XNOR2xp5_ASAP7_75t_R   g1024( .A (n1350), .B (n1355), .Y (y94) );
  INVx1_ASAP7_75t_R      g1025( .A (x222), .Y (n480) );
  NOR2xp33_ASAP7_75t_R   g1026( .A (n352), .B (n480), .Y (n1353) );
  NAND2xp33_ASAP7_75t_R  g1027( .A (x93), .B (x221), .Y (n1345) );
  NOR2xp33_ASAP7_75t_R   g1028( .A (x94), .B (x222), .Y (n1351) );
  NAND2xp33_ASAP7_75t_R  g1029( .A (n351), .B (n479), .Y (n1343) );
  OAI21xp33_ASAP7_75t_R  g1030( .A1 (n1335), .A2 (n1339), .B (n1343), .Y (n1349) );
  AOI21xp33_ASAP7_75t_R  g1031( .A1 (n1345), .B (n1351), .A2 (n1349), .Y (n1357) );
  NOR2xp33_ASAP7_75t_R   g1032( .A (n1353), .B (n1357), .Y (n1359) );
  INVx1_ASAP7_75t_R      g1033( .A (x95), .Y (n353) );
  XNOR2xp5_ASAP7_75t_R   g1034( .A (n353), .B (x223), .Y (n1364) );
  XNOR2xp5_ASAP7_75t_R   g1035( .A (n1359), .B (n1364), .Y (y95) );
  INVx1_ASAP7_75t_R      g1036( .A (x223), .Y (n481) );
  NOR2xp33_ASAP7_75t_R   g1037( .A (n353), .B (n481), .Y (n1362) );
  NAND2xp33_ASAP7_75t_R  g1038( .A (x94), .B (x222), .Y (n1354) );
  NOR2xp33_ASAP7_75t_R   g1039( .A (x95), .B (x223), .Y (n1360) );
  NAND2xp33_ASAP7_75t_R  g1040( .A (n352), .B (n480), .Y (n1352) );
  OAI21xp33_ASAP7_75t_R  g1041( .A1 (n1344), .A2 (n1348), .B (n1352), .Y (n1358) );
  AOI21xp33_ASAP7_75t_R  g1042( .A1 (n1354), .B (n1360), .A2 (n1358), .Y (n1366) );
  NOR2xp33_ASAP7_75t_R   g1043( .A (n1362), .B (n1366), .Y (n1368) );
  INVx1_ASAP7_75t_R      g1044( .A (x96), .Y (n354) );
  XNOR2xp5_ASAP7_75t_R   g1045( .A (n354), .B (x224), .Y (n1373) );
  XNOR2xp5_ASAP7_75t_R   g1046( .A (n1368), .B (n1373), .Y (y96) );
  INVx1_ASAP7_75t_R      g1047( .A (x224), .Y (n482) );
  NOR2xp33_ASAP7_75t_R   g1048( .A (n354), .B (n482), .Y (n1371) );
  NAND2xp33_ASAP7_75t_R  g1049( .A (x95), .B (x223), .Y (n1363) );
  NOR2xp33_ASAP7_75t_R   g1050( .A (x96), .B (x224), .Y (n1369) );
  NAND2xp33_ASAP7_75t_R  g1051( .A (n353), .B (n481), .Y (n1361) );
  OAI21xp33_ASAP7_75t_R  g1052( .A1 (n1353), .A2 (n1357), .B (n1361), .Y (n1367) );
  AOI21xp33_ASAP7_75t_R  g1053( .A1 (n1363), .B (n1369), .A2 (n1367), .Y (n1375) );
  NOR2xp33_ASAP7_75t_R   g1054( .A (n1371), .B (n1375), .Y (n1377) );
  INVx1_ASAP7_75t_R      g1055( .A (x97), .Y (n355) );
  XNOR2xp5_ASAP7_75t_R   g1056( .A (n355), .B (x225), .Y (n1382) );
  XNOR2xp5_ASAP7_75t_R   g1057( .A (n1377), .B (n1382), .Y (y97) );
  INVx1_ASAP7_75t_R      g1058( .A (x225), .Y (n483) );
  NOR2xp33_ASAP7_75t_R   g1059( .A (n355), .B (n483), .Y (n1380) );
  NAND2xp33_ASAP7_75t_R  g1060( .A (x96), .B (x224), .Y (n1372) );
  NOR2xp33_ASAP7_75t_R   g1061( .A (x97), .B (x225), .Y (n1378) );
  NAND2xp33_ASAP7_75t_R  g1062( .A (n354), .B (n482), .Y (n1370) );
  OAI21xp33_ASAP7_75t_R  g1063( .A1 (n1362), .A2 (n1366), .B (n1370), .Y (n1376) );
  AOI21xp33_ASAP7_75t_R  g1064( .A1 (n1372), .B (n1378), .A2 (n1376), .Y (n1384) );
  NOR2xp33_ASAP7_75t_R   g1065( .A (n1380), .B (n1384), .Y (n1386) );
  INVx1_ASAP7_75t_R      g1066( .A (x98), .Y (n356) );
  XNOR2xp5_ASAP7_75t_R   g1067( .A (n356), .B (x226), .Y (n1391) );
  XNOR2xp5_ASAP7_75t_R   g1068( .A (n1386), .B (n1391), .Y (y98) );
  INVx1_ASAP7_75t_R      g1069( .A (x226), .Y (n484) );
  NOR2xp33_ASAP7_75t_R   g1070( .A (n356), .B (n484), .Y (n1389) );
  NAND2xp33_ASAP7_75t_R  g1071( .A (x97), .B (x225), .Y (n1381) );
  NOR2xp33_ASAP7_75t_R   g1072( .A (x98), .B (x226), .Y (n1387) );
  NAND2xp33_ASAP7_75t_R  g1073( .A (n355), .B (n483), .Y (n1379) );
  OAI21xp33_ASAP7_75t_R  g1074( .A1 (n1371), .A2 (n1375), .B (n1379), .Y (n1385) );
  AOI21xp33_ASAP7_75t_R  g1075( .A1 (n1381), .B (n1387), .A2 (n1385), .Y (n1393) );
  NOR2xp33_ASAP7_75t_R   g1076( .A (n1389), .B (n1393), .Y (n1395) );
  INVx1_ASAP7_75t_R      g1077( .A (x99), .Y (n357) );
  XNOR2xp5_ASAP7_75t_R   g1078( .A (n357), .B (x227), .Y (n1400) );
  XNOR2xp5_ASAP7_75t_R   g1079( .A (n1395), .B (n1400), .Y (y99) );
  INVx1_ASAP7_75t_R      g1080( .A (x227), .Y (n485) );
  NOR2xp33_ASAP7_75t_R   g1081( .A (n357), .B (n485), .Y (n1398) );
  NAND2xp33_ASAP7_75t_R  g1082( .A (x98), .B (x226), .Y (n1390) );
  NOR2xp33_ASAP7_75t_R   g1083( .A (x99), .B (x227), .Y (n1396) );
  NAND2xp33_ASAP7_75t_R  g1084( .A (n356), .B (n484), .Y (n1388) );
  OAI21xp33_ASAP7_75t_R  g1085( .A1 (n1380), .A2 (n1384), .B (n1388), .Y (n1394) );
  AOI21xp33_ASAP7_75t_R  g1086( .A1 (n1390), .B (n1396), .A2 (n1394), .Y (n1402) );
  NOR2xp33_ASAP7_75t_R   g1087( .A (n1398), .B (n1402), .Y (n1404) );
  INVx1_ASAP7_75t_R      g1088( .A (x100), .Y (n358) );
  XNOR2xp5_ASAP7_75t_R   g1089( .A (n358), .B (x228), .Y (n1409) );
  XNOR2xp5_ASAP7_75t_R   g1090( .A (n1404), .B (n1409), .Y (y100) );
  INVx1_ASAP7_75t_R      g1091( .A (x228), .Y (n486) );
  NOR2xp33_ASAP7_75t_R   g1092( .A (n358), .B (n486), .Y (n1407) );
  NAND2xp33_ASAP7_75t_R  g1093( .A (x99), .B (x227), .Y (n1399) );
  NOR2xp33_ASAP7_75t_R   g1094( .A (x100), .B (x228), .Y (n1405) );
  NAND2xp33_ASAP7_75t_R  g1095( .A (n357), .B (n485), .Y (n1397) );
  OAI21xp33_ASAP7_75t_R  g1096( .A1 (n1389), .A2 (n1393), .B (n1397), .Y (n1403) );
  AOI21xp33_ASAP7_75t_R  g1097( .A1 (n1399), .B (n1405), .A2 (n1403), .Y (n1411) );
  NOR2xp33_ASAP7_75t_R   g1098( .A (n1407), .B (n1411), .Y (n1413) );
  INVx1_ASAP7_75t_R      g1099( .A (x101), .Y (n359) );
  XNOR2xp5_ASAP7_75t_R   g1100( .A (n359), .B (x229), .Y (n1418) );
  XNOR2xp5_ASAP7_75t_R   g1101( .A (n1413), .B (n1418), .Y (y101) );
  INVx1_ASAP7_75t_R      g1102( .A (x229), .Y (n487) );
  NOR2xp33_ASAP7_75t_R   g1103( .A (n359), .B (n487), .Y (n1416) );
  NAND2xp33_ASAP7_75t_R  g1104( .A (x100), .B (x228), .Y (n1408) );
  NOR2xp33_ASAP7_75t_R   g1105( .A (x101), .B (x229), .Y (n1414) );
  NAND2xp33_ASAP7_75t_R  g1106( .A (n358), .B (n486), .Y (n1406) );
  OAI21xp33_ASAP7_75t_R  g1107( .A1 (n1398), .A2 (n1402), .B (n1406), .Y (n1412) );
  AOI21xp33_ASAP7_75t_R  g1108( .A1 (n1408), .B (n1414), .A2 (n1412), .Y (n1420) );
  NOR2xp33_ASAP7_75t_R   g1109( .A (n1416), .B (n1420), .Y (n1422) );
  INVx1_ASAP7_75t_R      g1110( .A (x102), .Y (n360) );
  XNOR2xp5_ASAP7_75t_R   g1111( .A (n360), .B (x230), .Y (n1427) );
  XNOR2xp5_ASAP7_75t_R   g1112( .A (n1422), .B (n1427), .Y (y102) );
  INVx1_ASAP7_75t_R      g1113( .A (x230), .Y (n488) );
  NOR2xp33_ASAP7_75t_R   g1114( .A (n360), .B (n488), .Y (n1425) );
  NAND2xp33_ASAP7_75t_R  g1115( .A (x101), .B (x229), .Y (n1417) );
  NOR2xp33_ASAP7_75t_R   g1116( .A (x102), .B (x230), .Y (n1423) );
  NAND2xp33_ASAP7_75t_R  g1117( .A (n359), .B (n487), .Y (n1415) );
  OAI21xp33_ASAP7_75t_R  g1118( .A1 (n1407), .A2 (n1411), .B (n1415), .Y (n1421) );
  AOI21xp33_ASAP7_75t_R  g1119( .A1 (n1417), .B (n1423), .A2 (n1421), .Y (n1429) );
  NOR2xp33_ASAP7_75t_R   g1120( .A (n1425), .B (n1429), .Y (n1431) );
  INVx1_ASAP7_75t_R      g1121( .A (x103), .Y (n361) );
  XNOR2xp5_ASAP7_75t_R   g1122( .A (n361), .B (x231), .Y (n1436) );
  XNOR2xp5_ASAP7_75t_R   g1123( .A (n1431), .B (n1436), .Y (y103) );
  INVx1_ASAP7_75t_R      g1124( .A (x231), .Y (n489) );
  NOR2xp33_ASAP7_75t_R   g1125( .A (n361), .B (n489), .Y (n1434) );
  NAND2xp33_ASAP7_75t_R  g1126( .A (x102), .B (x230), .Y (n1426) );
  NOR2xp33_ASAP7_75t_R   g1127( .A (x103), .B (x231), .Y (n1432) );
  NAND2xp33_ASAP7_75t_R  g1128( .A (n360), .B (n488), .Y (n1424) );
  OAI21xp33_ASAP7_75t_R  g1129( .A1 (n1416), .A2 (n1420), .B (n1424), .Y (n1430) );
  AOI21xp33_ASAP7_75t_R  g1130( .A1 (n1426), .B (n1432), .A2 (n1430), .Y (n1438) );
  NOR2xp33_ASAP7_75t_R   g1131( .A (n1434), .B (n1438), .Y (n1440) );
  INVx1_ASAP7_75t_R      g1132( .A (x104), .Y (n362) );
  XNOR2xp5_ASAP7_75t_R   g1133( .A (n362), .B (x232), .Y (n1445) );
  XNOR2xp5_ASAP7_75t_R   g1134( .A (n1440), .B (n1445), .Y (y104) );
  INVx1_ASAP7_75t_R      g1135( .A (x232), .Y (n490) );
  NOR2xp33_ASAP7_75t_R   g1136( .A (n362), .B (n490), .Y (n1443) );
  NAND2xp33_ASAP7_75t_R  g1137( .A (x103), .B (x231), .Y (n1435) );
  NOR2xp33_ASAP7_75t_R   g1138( .A (x104), .B (x232), .Y (n1441) );
  NAND2xp33_ASAP7_75t_R  g1139( .A (n361), .B (n489), .Y (n1433) );
  OAI21xp33_ASAP7_75t_R  g1140( .A1 (n1425), .A2 (n1429), .B (n1433), .Y (n1439) );
  AOI21xp33_ASAP7_75t_R  g1141( .A1 (n1435), .B (n1441), .A2 (n1439), .Y (n1447) );
  NOR2xp33_ASAP7_75t_R   g1142( .A (n1443), .B (n1447), .Y (n1449) );
  INVx1_ASAP7_75t_R      g1143( .A (x105), .Y (n363) );
  XNOR2xp5_ASAP7_75t_R   g1144( .A (n363), .B (x233), .Y (n1454) );
  XNOR2xp5_ASAP7_75t_R   g1145( .A (n1449), .B (n1454), .Y (y105) );
  INVx1_ASAP7_75t_R      g1146( .A (x233), .Y (n491) );
  NOR2xp33_ASAP7_75t_R   g1147( .A (n363), .B (n491), .Y (n1452) );
  NAND2xp33_ASAP7_75t_R  g1148( .A (x104), .B (x232), .Y (n1444) );
  NOR2xp33_ASAP7_75t_R   g1149( .A (x105), .B (x233), .Y (n1450) );
  NAND2xp33_ASAP7_75t_R  g1150( .A (n362), .B (n490), .Y (n1442) );
  OAI21xp33_ASAP7_75t_R  g1151( .A1 (n1434), .A2 (n1438), .B (n1442), .Y (n1448) );
  AOI21xp33_ASAP7_75t_R  g1152( .A1 (n1444), .B (n1450), .A2 (n1448), .Y (n1456) );
  NOR2xp33_ASAP7_75t_R   g1153( .A (n1452), .B (n1456), .Y (n1458) );
  INVx1_ASAP7_75t_R      g1154( .A (x106), .Y (n364) );
  XNOR2xp5_ASAP7_75t_R   g1155( .A (n364), .B (x234), .Y (n1463) );
  XNOR2xp5_ASAP7_75t_R   g1156( .A (n1458), .B (n1463), .Y (y106) );
  INVx1_ASAP7_75t_R      g1157( .A (x234), .Y (n492) );
  NOR2xp33_ASAP7_75t_R   g1158( .A (n364), .B (n492), .Y (n1461) );
  NAND2xp33_ASAP7_75t_R  g1159( .A (x105), .B (x233), .Y (n1453) );
  NOR2xp33_ASAP7_75t_R   g1160( .A (x106), .B (x234), .Y (n1459) );
  NAND2xp33_ASAP7_75t_R  g1161( .A (n363), .B (n491), .Y (n1451) );
  OAI21xp33_ASAP7_75t_R  g1162( .A1 (n1443), .A2 (n1447), .B (n1451), .Y (n1457) );
  AOI21xp33_ASAP7_75t_R  g1163( .A1 (n1453), .B (n1459), .A2 (n1457), .Y (n1465) );
  NOR2xp33_ASAP7_75t_R   g1164( .A (n1461), .B (n1465), .Y (n1467) );
  INVx1_ASAP7_75t_R      g1165( .A (x107), .Y (n365) );
  XNOR2xp5_ASAP7_75t_R   g1166( .A (n365), .B (x235), .Y (n1472) );
  XNOR2xp5_ASAP7_75t_R   g1167( .A (n1467), .B (n1472), .Y (y107) );
  INVx1_ASAP7_75t_R      g1168( .A (x235), .Y (n493) );
  NOR2xp33_ASAP7_75t_R   g1169( .A (n365), .B (n493), .Y (n1470) );
  NAND2xp33_ASAP7_75t_R  g1170( .A (x106), .B (x234), .Y (n1462) );
  NOR2xp33_ASAP7_75t_R   g1171( .A (x107), .B (x235), .Y (n1468) );
  NAND2xp33_ASAP7_75t_R  g1172( .A (n364), .B (n492), .Y (n1460) );
  OAI21xp33_ASAP7_75t_R  g1173( .A1 (n1452), .A2 (n1456), .B (n1460), .Y (n1466) );
  AOI21xp33_ASAP7_75t_R  g1174( .A1 (n1462), .B (n1468), .A2 (n1466), .Y (n1474) );
  NOR2xp33_ASAP7_75t_R   g1175( .A (n1470), .B (n1474), .Y (n1476) );
  INVx1_ASAP7_75t_R      g1176( .A (x108), .Y (n366) );
  XNOR2xp5_ASAP7_75t_R   g1177( .A (n366), .B (x236), .Y (n1481) );
  XNOR2xp5_ASAP7_75t_R   g1178( .A (n1476), .B (n1481), .Y (y108) );
  INVx1_ASAP7_75t_R      g1179( .A (x236), .Y (n494) );
  NOR2xp33_ASAP7_75t_R   g1180( .A (n366), .B (n494), .Y (n1479) );
  NAND2xp33_ASAP7_75t_R  g1181( .A (x107), .B (x235), .Y (n1471) );
  NOR2xp33_ASAP7_75t_R   g1182( .A (x108), .B (x236), .Y (n1477) );
  NAND2xp33_ASAP7_75t_R  g1183( .A (n365), .B (n493), .Y (n1469) );
  OAI21xp33_ASAP7_75t_R  g1184( .A1 (n1461), .A2 (n1465), .B (n1469), .Y (n1475) );
  AOI21xp33_ASAP7_75t_R  g1185( .A1 (n1471), .B (n1477), .A2 (n1475), .Y (n1483) );
  NOR2xp33_ASAP7_75t_R   g1186( .A (n1479), .B (n1483), .Y (n1485) );
  INVx1_ASAP7_75t_R      g1187( .A (x109), .Y (n367) );
  XNOR2xp5_ASAP7_75t_R   g1188( .A (n367), .B (x237), .Y (n1490) );
  XNOR2xp5_ASAP7_75t_R   g1189( .A (n1485), .B (n1490), .Y (y109) );
  INVx1_ASAP7_75t_R      g1190( .A (x237), .Y (n495) );
  NOR2xp33_ASAP7_75t_R   g1191( .A (n367), .B (n495), .Y (n1488) );
  NAND2xp33_ASAP7_75t_R  g1192( .A (x108), .B (x236), .Y (n1480) );
  NOR2xp33_ASAP7_75t_R   g1193( .A (x109), .B (x237), .Y (n1486) );
  NAND2xp33_ASAP7_75t_R  g1194( .A (n366), .B (n494), .Y (n1478) );
  OAI21xp33_ASAP7_75t_R  g1195( .A1 (n1470), .A2 (n1474), .B (n1478), .Y (n1484) );
  AOI21xp33_ASAP7_75t_R  g1196( .A1 (n1480), .B (n1486), .A2 (n1484), .Y (n1492) );
  NOR2xp33_ASAP7_75t_R   g1197( .A (n1488), .B (n1492), .Y (n1494) );
  INVx1_ASAP7_75t_R      g1198( .A (x110), .Y (n368) );
  XNOR2xp5_ASAP7_75t_R   g1199( .A (n368), .B (x238), .Y (n1499) );
  XNOR2xp5_ASAP7_75t_R   g1200( .A (n1494), .B (n1499), .Y (y110) );
  INVx1_ASAP7_75t_R      g1201( .A (x238), .Y (n496) );
  NOR2xp33_ASAP7_75t_R   g1202( .A (n368), .B (n496), .Y (n1497) );
  NAND2xp33_ASAP7_75t_R  g1203( .A (x109), .B (x237), .Y (n1489) );
  NOR2xp33_ASAP7_75t_R   g1204( .A (x110), .B (x238), .Y (n1495) );
  NAND2xp33_ASAP7_75t_R  g1205( .A (n367), .B (n495), .Y (n1487) );
  OAI21xp33_ASAP7_75t_R  g1206( .A1 (n1479), .A2 (n1483), .B (n1487), .Y (n1493) );
  AOI21xp33_ASAP7_75t_R  g1207( .A1 (n1489), .B (n1495), .A2 (n1493), .Y (n1501) );
  NOR2xp33_ASAP7_75t_R   g1208( .A (n1497), .B (n1501), .Y (n1503) );
  INVx1_ASAP7_75t_R      g1209( .A (x111), .Y (n369) );
  XNOR2xp5_ASAP7_75t_R   g1210( .A (n369), .B (x239), .Y (n1508) );
  XNOR2xp5_ASAP7_75t_R   g1211( .A (n1503), .B (n1508), .Y (y111) );
  INVx1_ASAP7_75t_R      g1212( .A (x239), .Y (n497) );
  NOR2xp33_ASAP7_75t_R   g1213( .A (n369), .B (n497), .Y (n1506) );
  NAND2xp33_ASAP7_75t_R  g1214( .A (x110), .B (x238), .Y (n1498) );
  NOR2xp33_ASAP7_75t_R   g1215( .A (x111), .B (x239), .Y (n1504) );
  NAND2xp33_ASAP7_75t_R  g1216( .A (n368), .B (n496), .Y (n1496) );
  OAI21xp33_ASAP7_75t_R  g1217( .A1 (n1488), .A2 (n1492), .B (n1496), .Y (n1502) );
  AOI21xp33_ASAP7_75t_R  g1218( .A1 (n1498), .B (n1504), .A2 (n1502), .Y (n1510) );
  NOR2xp33_ASAP7_75t_R   g1219( .A (n1506), .B (n1510), .Y (n1512) );
  INVx1_ASAP7_75t_R      g1220( .A (x112), .Y (n370) );
  XNOR2xp5_ASAP7_75t_R   g1221( .A (n370), .B (x240), .Y (n1517) );
  XNOR2xp5_ASAP7_75t_R   g1222( .A (n1512), .B (n1517), .Y (y112) );
  INVx1_ASAP7_75t_R      g1223( .A (x240), .Y (n498) );
  NOR2xp33_ASAP7_75t_R   g1224( .A (n370), .B (n498), .Y (n1515) );
  NAND2xp33_ASAP7_75t_R  g1225( .A (x111), .B (x239), .Y (n1507) );
  NOR2xp33_ASAP7_75t_R   g1226( .A (x112), .B (x240), .Y (n1513) );
  NAND2xp33_ASAP7_75t_R  g1227( .A (n369), .B (n497), .Y (n1505) );
  OAI21xp33_ASAP7_75t_R  g1228( .A1 (n1497), .A2 (n1501), .B (n1505), .Y (n1511) );
  AOI21xp33_ASAP7_75t_R  g1229( .A1 (n1507), .B (n1513), .A2 (n1511), .Y (n1519) );
  NOR2xp33_ASAP7_75t_R   g1230( .A (n1515), .B (n1519), .Y (n1521) );
  INVx1_ASAP7_75t_R      g1231( .A (x113), .Y (n371) );
  XNOR2xp5_ASAP7_75t_R   g1232( .A (n371), .B (x241), .Y (n1526) );
  XNOR2xp5_ASAP7_75t_R   g1233( .A (n1521), .B (n1526), .Y (y113) );
  INVx1_ASAP7_75t_R      g1234( .A (x241), .Y (n499) );
  NOR2xp33_ASAP7_75t_R   g1235( .A (n371), .B (n499), .Y (n1524) );
  NAND2xp33_ASAP7_75t_R  g1236( .A (x112), .B (x240), .Y (n1516) );
  NOR2xp33_ASAP7_75t_R   g1237( .A (x113), .B (x241), .Y (n1522) );
  NAND2xp33_ASAP7_75t_R  g1238( .A (n370), .B (n498), .Y (n1514) );
  OAI21xp33_ASAP7_75t_R  g1239( .A1 (n1506), .A2 (n1510), .B (n1514), .Y (n1520) );
  AOI21xp33_ASAP7_75t_R  g1240( .A1 (n1516), .B (n1522), .A2 (n1520), .Y (n1528) );
  NOR2xp33_ASAP7_75t_R   g1241( .A (n1524), .B (n1528), .Y (n1530) );
  INVx1_ASAP7_75t_R      g1242( .A (x114), .Y (n372) );
  XNOR2xp5_ASAP7_75t_R   g1243( .A (n372), .B (x242), .Y (n1535) );
  XNOR2xp5_ASAP7_75t_R   g1244( .A (n1530), .B (n1535), .Y (y114) );
  INVx1_ASAP7_75t_R      g1245( .A (x242), .Y (n500) );
  NOR2xp33_ASAP7_75t_R   g1246( .A (n372), .B (n500), .Y (n1533) );
  NAND2xp33_ASAP7_75t_R  g1247( .A (x113), .B (x241), .Y (n1525) );
  NOR2xp33_ASAP7_75t_R   g1248( .A (x114), .B (x242), .Y (n1531) );
  NAND2xp33_ASAP7_75t_R  g1249( .A (n371), .B (n499), .Y (n1523) );
  OAI21xp33_ASAP7_75t_R  g1250( .A1 (n1515), .A2 (n1519), .B (n1523), .Y (n1529) );
  AOI21xp33_ASAP7_75t_R  g1251( .A1 (n1525), .B (n1531), .A2 (n1529), .Y (n1537) );
  NOR2xp33_ASAP7_75t_R   g1252( .A (n1533), .B (n1537), .Y (n1539) );
  INVx1_ASAP7_75t_R      g1253( .A (x115), .Y (n373) );
  XNOR2xp5_ASAP7_75t_R   g1254( .A (n373), .B (x243), .Y (n1544) );
  XNOR2xp5_ASAP7_75t_R   g1255( .A (n1539), .B (n1544), .Y (y115) );
  INVx1_ASAP7_75t_R      g1256( .A (x243), .Y (n501) );
  NOR2xp33_ASAP7_75t_R   g1257( .A (n373), .B (n501), .Y (n1542) );
  NAND2xp33_ASAP7_75t_R  g1258( .A (x114), .B (x242), .Y (n1534) );
  NOR2xp33_ASAP7_75t_R   g1259( .A (x115), .B (x243), .Y (n1540) );
  NAND2xp33_ASAP7_75t_R  g1260( .A (n372), .B (n500), .Y (n1532) );
  OAI21xp33_ASAP7_75t_R  g1261( .A1 (n1524), .A2 (n1528), .B (n1532), .Y (n1538) );
  AOI21xp33_ASAP7_75t_R  g1262( .A1 (n1534), .B (n1540), .A2 (n1538), .Y (n1546) );
  NOR2xp33_ASAP7_75t_R   g1263( .A (n1542), .B (n1546), .Y (n1548) );
  INVx1_ASAP7_75t_R      g1264( .A (x116), .Y (n374) );
  XNOR2xp5_ASAP7_75t_R   g1265( .A (n374), .B (x244), .Y (n1553) );
  XNOR2xp5_ASAP7_75t_R   g1266( .A (n1548), .B (n1553), .Y (y116) );
  INVx1_ASAP7_75t_R      g1267( .A (x244), .Y (n502) );
  NOR2xp33_ASAP7_75t_R   g1268( .A (n374), .B (n502), .Y (n1551) );
  NAND2xp33_ASAP7_75t_R  g1269( .A (x115), .B (x243), .Y (n1543) );
  NOR2xp33_ASAP7_75t_R   g1270( .A (x116), .B (x244), .Y (n1549) );
  NAND2xp33_ASAP7_75t_R  g1271( .A (n373), .B (n501), .Y (n1541) );
  OAI21xp33_ASAP7_75t_R  g1272( .A1 (n1533), .A2 (n1537), .B (n1541), .Y (n1547) );
  AOI21xp33_ASAP7_75t_R  g1273( .A1 (n1543), .B (n1549), .A2 (n1547), .Y (n1555) );
  NOR2xp33_ASAP7_75t_R   g1274( .A (n1551), .B (n1555), .Y (n1557) );
  INVx1_ASAP7_75t_R      g1275( .A (x117), .Y (n375) );
  XNOR2xp5_ASAP7_75t_R   g1276( .A (n375), .B (x245), .Y (n1562) );
  XNOR2xp5_ASAP7_75t_R   g1277( .A (n1557), .B (n1562), .Y (y117) );
  INVx1_ASAP7_75t_R      g1278( .A (x245), .Y (n503) );
  NOR2xp33_ASAP7_75t_R   g1279( .A (n375), .B (n503), .Y (n1560) );
  NAND2xp33_ASAP7_75t_R  g1280( .A (x116), .B (x244), .Y (n1552) );
  NOR2xp33_ASAP7_75t_R   g1281( .A (x117), .B (x245), .Y (n1558) );
  NAND2xp33_ASAP7_75t_R  g1282( .A (n374), .B (n502), .Y (n1550) );
  OAI21xp33_ASAP7_75t_R  g1283( .A1 (n1542), .A2 (n1546), .B (n1550), .Y (n1556) );
  AOI21xp33_ASAP7_75t_R  g1284( .A1 (n1552), .B (n1558), .A2 (n1556), .Y (n1564) );
  NOR2xp33_ASAP7_75t_R   g1285( .A (n1560), .B (n1564), .Y (n1566) );
  INVx1_ASAP7_75t_R      g1286( .A (x118), .Y (n376) );
  XNOR2xp5_ASAP7_75t_R   g1287( .A (n376), .B (x246), .Y (n1571) );
  XNOR2xp5_ASAP7_75t_R   g1288( .A (n1566), .B (n1571), .Y (y118) );
  INVx1_ASAP7_75t_R      g1289( .A (x246), .Y (n504) );
  NOR2xp33_ASAP7_75t_R   g1290( .A (n376), .B (n504), .Y (n1569) );
  NAND2xp33_ASAP7_75t_R  g1291( .A (x117), .B (x245), .Y (n1561) );
  NOR2xp33_ASAP7_75t_R   g1292( .A (x118), .B (x246), .Y (n1567) );
  NAND2xp33_ASAP7_75t_R  g1293( .A (n375), .B (n503), .Y (n1559) );
  OAI21xp33_ASAP7_75t_R  g1294( .A1 (n1551), .A2 (n1555), .B (n1559), .Y (n1565) );
  AOI21xp33_ASAP7_75t_R  g1295( .A1 (n1561), .B (n1567), .A2 (n1565), .Y (n1573) );
  NOR2xp33_ASAP7_75t_R   g1296( .A (n1569), .B (n1573), .Y (n1575) );
  INVx1_ASAP7_75t_R      g1297( .A (x119), .Y (n377) );
  XNOR2xp5_ASAP7_75t_R   g1298( .A (n377), .B (x247), .Y (n1580) );
  XNOR2xp5_ASAP7_75t_R   g1299( .A (n1575), .B (n1580), .Y (y119) );
  INVx1_ASAP7_75t_R      g1300( .A (x247), .Y (n505) );
  NOR2xp33_ASAP7_75t_R   g1301( .A (n377), .B (n505), .Y (n1578) );
  NAND2xp33_ASAP7_75t_R  g1302( .A (x118), .B (x246), .Y (n1570) );
  NOR2xp33_ASAP7_75t_R   g1303( .A (x119), .B (x247), .Y (n1576) );
  NAND2xp33_ASAP7_75t_R  g1304( .A (n376), .B (n504), .Y (n1568) );
  OAI21xp33_ASAP7_75t_R  g1305( .A1 (n1560), .A2 (n1564), .B (n1568), .Y (n1574) );
  AOI21xp33_ASAP7_75t_R  g1306( .A1 (n1570), .B (n1576), .A2 (n1574), .Y (n1582) );
  NOR2xp33_ASAP7_75t_R   g1307( .A (n1578), .B (n1582), .Y (n1584) );
  INVx1_ASAP7_75t_R      g1308( .A (x120), .Y (n378) );
  XNOR2xp5_ASAP7_75t_R   g1309( .A (n378), .B (x248), .Y (n1589) );
  XNOR2xp5_ASAP7_75t_R   g1310( .A (n1584), .B (n1589), .Y (y120) );
  INVx1_ASAP7_75t_R      g1311( .A (x248), .Y (n506) );
  NOR2xp33_ASAP7_75t_R   g1312( .A (n378), .B (n506), .Y (n1587) );
  NAND2xp33_ASAP7_75t_R  g1313( .A (x119), .B (x247), .Y (n1579) );
  NOR2xp33_ASAP7_75t_R   g1314( .A (x120), .B (x248), .Y (n1585) );
  NAND2xp33_ASAP7_75t_R  g1315( .A (n377), .B (n505), .Y (n1577) );
  OAI21xp33_ASAP7_75t_R  g1316( .A1 (n1569), .A2 (n1573), .B (n1577), .Y (n1583) );
  AOI21xp33_ASAP7_75t_R  g1317( .A1 (n1579), .B (n1585), .A2 (n1583), .Y (n1591) );
  NOR2xp33_ASAP7_75t_R   g1318( .A (n1587), .B (n1591), .Y (n1593) );
  INVx1_ASAP7_75t_R      g1319( .A (x121), .Y (n379) );
  XNOR2xp5_ASAP7_75t_R   g1320( .A (n379), .B (x249), .Y (n1598) );
  XNOR2xp5_ASAP7_75t_R   g1321( .A (n1593), .B (n1598), .Y (y121) );
  INVx1_ASAP7_75t_R      g1322( .A (x249), .Y (n507) );
  NOR2xp33_ASAP7_75t_R   g1323( .A (n379), .B (n507), .Y (n1596) );
  NAND2xp33_ASAP7_75t_R  g1324( .A (x120), .B (x248), .Y (n1588) );
  NOR2xp33_ASAP7_75t_R   g1325( .A (x121), .B (x249), .Y (n1594) );
  NAND2xp33_ASAP7_75t_R  g1326( .A (n378), .B (n506), .Y (n1586) );
  OAI21xp33_ASAP7_75t_R  g1327( .A1 (n1578), .A2 (n1582), .B (n1586), .Y (n1592) );
  AOI21xp33_ASAP7_75t_R  g1328( .A1 (n1588), .B (n1594), .A2 (n1592), .Y (n1600) );
  NOR2xp33_ASAP7_75t_R   g1329( .A (n1596), .B (n1600), .Y (n1602) );
  INVx1_ASAP7_75t_R      g1330( .A (x122), .Y (n380) );
  XNOR2xp5_ASAP7_75t_R   g1331( .A (n380), .B (x250), .Y (n1607) );
  XNOR2xp5_ASAP7_75t_R   g1332( .A (n1602), .B (n1607), .Y (y122) );
  INVx1_ASAP7_75t_R      g1333( .A (x250), .Y (n508) );
  NOR2xp33_ASAP7_75t_R   g1334( .A (n380), .B (n508), .Y (n1605) );
  NAND2xp33_ASAP7_75t_R  g1335( .A (x121), .B (x249), .Y (n1597) );
  NOR2xp33_ASAP7_75t_R   g1336( .A (x122), .B (x250), .Y (n1603) );
  NAND2xp33_ASAP7_75t_R  g1337( .A (n379), .B (n507), .Y (n1595) );
  OAI21xp33_ASAP7_75t_R  g1338( .A1 (n1587), .A2 (n1591), .B (n1595), .Y (n1601) );
  AOI21xp33_ASAP7_75t_R  g1339( .A1 (n1597), .B (n1603), .A2 (n1601), .Y (n1609) );
  NOR2xp33_ASAP7_75t_R   g1340( .A (n1605), .B (n1609), .Y (n1611) );
  INVx1_ASAP7_75t_R      g1341( .A (x123), .Y (n381) );
  XNOR2xp5_ASAP7_75t_R   g1342( .A (n381), .B (x251), .Y (n1616) );
  XNOR2xp5_ASAP7_75t_R   g1343( .A (n1611), .B (n1616), .Y (y123) );
  INVx1_ASAP7_75t_R      g1344( .A (x251), .Y (n509) );
  NOR2xp33_ASAP7_75t_R   g1345( .A (n381), .B (n509), .Y (n1614) );
  NAND2xp33_ASAP7_75t_R  g1346( .A (x122), .B (x250), .Y (n1606) );
  NOR2xp33_ASAP7_75t_R   g1347( .A (x123), .B (x251), .Y (n1612) );
  NAND2xp33_ASAP7_75t_R  g1348( .A (n380), .B (n508), .Y (n1604) );
  OAI21xp33_ASAP7_75t_R  g1349( .A1 (n1596), .A2 (n1600), .B (n1604), .Y (n1610) );
  AOI21xp33_ASAP7_75t_R  g1350( .A1 (n1606), .B (n1612), .A2 (n1610), .Y (n1618) );
  NOR2xp33_ASAP7_75t_R   g1351( .A (n1614), .B (n1618), .Y (n1620) );
  INVx1_ASAP7_75t_R      g1352( .A (x124), .Y (n382) );
  XNOR2xp5_ASAP7_75t_R   g1353( .A (n382), .B (x252), .Y (n1625) );
  XNOR2xp5_ASAP7_75t_R   g1354( .A (n1620), .B (n1625), .Y (y124) );
  INVx1_ASAP7_75t_R      g1355( .A (x252), .Y (n510) );
  NOR2xp33_ASAP7_75t_R   g1356( .A (n382), .B (n510), .Y (n1623) );
  NAND2xp33_ASAP7_75t_R  g1357( .A (x123), .B (x251), .Y (n1615) );
  NOR2xp33_ASAP7_75t_R   g1358( .A (x124), .B (x252), .Y (n1621) );
  NAND2xp33_ASAP7_75t_R  g1359( .A (n381), .B (n509), .Y (n1613) );
  OAI21xp33_ASAP7_75t_R  g1360( .A1 (n1605), .A2 (n1609), .B (n1613), .Y (n1619) );
  AOI21xp33_ASAP7_75t_R  g1361( .A1 (n1615), .B (n1621), .A2 (n1619), .Y (n1627) );
  NOR2xp33_ASAP7_75t_R   g1362( .A (n1623), .B (n1627), .Y (n1629) );
  INVx1_ASAP7_75t_R      g1363( .A (x125), .Y (n383) );
  XNOR2xp5_ASAP7_75t_R   g1364( .A (n383), .B (x253), .Y (n1634) );
  XNOR2xp5_ASAP7_75t_R   g1365( .A (n1629), .B (n1634), .Y (y125) );
  INVx1_ASAP7_75t_R      g1366( .A (x253), .Y (n511) );
  NOR2xp33_ASAP7_75t_R   g1367( .A (n383), .B (n511), .Y (n1632) );
  NAND2xp33_ASAP7_75t_R  g1368( .A (x124), .B (x252), .Y (n1624) );
  NOR2xp33_ASAP7_75t_R   g1369( .A (x125), .B (x253), .Y (n1630) );
  NAND2xp33_ASAP7_75t_R  g1370( .A (n382), .B (n510), .Y (n1622) );
  OAI21xp33_ASAP7_75t_R  g1371( .A1 (n1614), .A2 (n1618), .B (n1622), .Y (n1628) );
  AOI21xp33_ASAP7_75t_R  g1372( .A1 (n1624), .B (n1630), .A2 (n1628), .Y (n1636) );
  NOR2xp33_ASAP7_75t_R   g1373( .A (n1632), .B (n1636), .Y (n1638) );
  INVx1_ASAP7_75t_R      g1374( .A (x126), .Y (n384) );
  XNOR2xp5_ASAP7_75t_R   g1375( .A (n384), .B (x254), .Y (n1641) );
  XNOR2xp5_ASAP7_75t_R   g1376( .A (n1638), .B (n1641), .Y (y126) );
  INVx1_ASAP7_75t_R      g1377( .A (x254), .Y (n512) );
  NOR2xp33_ASAP7_75t_R   g1378( .A (n384), .B (n512), .Y (n1640) );
  NAND2xp33_ASAP7_75t_R  g1379( .A (x125), .B (x253), .Y (n1633) );
  NOR2xp33_ASAP7_75t_R   g1380( .A (x126), .B (x254), .Y (n1639) );
  NAND2xp33_ASAP7_75t_R  g1381( .A (n383), .B (n511), .Y (n1631) );
  OAI21xp33_ASAP7_75t_R  g1382( .A1 (n1623), .A2 (n1627), .B (n1631), .Y (n1637) );
  AOI21xp33_ASAP7_75t_R  g1383( .A1 (n1633), .B (n1639), .A2 (n1637), .Y (n1643) );
  NOR2xp33_ASAP7_75t_R   g1384( .A (n1640), .B (n1643), .Y (n1644) );
  INVx1_ASAP7_75t_R      g1385( .A (x127), .Y (n385) );
  XNOR2xp5_ASAP7_75t_R   g1386( .A (n385), .B (x255), .Y (n1647) );
  XNOR2xp5_ASAP7_75t_R   g1387( .A (n1644), .B (n1647), .Y (y127) );
  NAND2xp33_ASAP7_75t_R  g1388( .A (x127), .B (x255), .Y (n1646) );
  INVx1_ASAP7_75t_R      g1389( .A (x255), .Y (n513) );
  NAND2xp33_ASAP7_75t_R  g1390( .A (n385), .B (n513), .Y (n1645) );
  OAI21xp33_ASAP7_75t_R  g1391( .A1 (n1640), .A2 (n1643), .B (n1645), .Y (n1649) );
  NAND2xp33_ASAP7_75t_R  g1392( .A (n1646), .B (n1649), .Y (y128) );
endmodule
